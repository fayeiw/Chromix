magic
tech sky130A
magscale 1 2
timestamp 1746053276
<< obsli1 >>
rect 1104 2159 22264 22865
<< obsm1 >>
rect 14 2128 22264 22896
<< metal2 >>
rect 1306 24752 1362 25552
rect 10322 24752 10378 25552
rect 19338 24752 19394 25552
rect 18 0 74 800
rect 8390 0 8446 800
rect 17406 0 17462 800
<< obsm2 >>
rect 20 24696 1250 24752
rect 1418 24696 10266 24752
rect 10434 24696 19282 24752
rect 19450 24696 22246 24752
rect 20 856 22246 24696
rect 130 734 8334 856
rect 8502 734 17350 856
rect 17518 734 22246 856
<< metal3 >>
rect 22608 21088 23408 21208
rect 0 18368 800 18488
rect 22608 11568 23408 11688
rect 0 8848 800 8968
rect 22608 2048 23408 2168
<< obsm3 >>
rect 800 21288 22608 22881
rect 800 21008 22528 21288
rect 800 18568 22608 21008
rect 880 18288 22608 18568
rect 800 11768 22608 18288
rect 800 11488 22528 11768
rect 800 9048 22608 11488
rect 880 8768 22608 9048
rect 800 2248 22608 8768
rect 800 2075 22528 2248
<< metal4 >>
rect 3589 2128 3909 22896
rect 4249 2128 4569 22896
rect 8879 2128 9199 22896
rect 9539 2128 9859 22896
rect 14169 2128 14489 22896
rect 14829 2128 15149 22896
rect 19459 2128 19779 22896
rect 20119 2128 20439 22896
<< metal5 >>
rect 1056 20764 22312 21084
rect 1056 20104 22312 20424
rect 1056 15596 22312 15916
rect 1056 14936 22312 15256
rect 1056 10428 22312 10748
rect 1056 9768 22312 10088
rect 1056 5260 22312 5580
rect 1056 4600 22312 4920
<< labels >>
rlabel metal4 s 4249 2128 4569 22896 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 9539 2128 9859 22896 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 14829 2128 15149 22896 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 20119 2128 20439 22896 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5260 22312 5580 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 10428 22312 10748 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 15596 22312 15916 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 20764 22312 21084 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3589 2128 3909 22896 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 8879 2128 9199 22896 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 14169 2128 14489 22896 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19459 2128 19779 22896 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4600 22312 4920 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 9768 22312 10088 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 14936 22312 15256 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 20104 22312 20424 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 18368 800 18488 6 clk
port 3 nsew signal input
rlabel metal3 s 22608 2048 23408 2168 6 enc0_a
port 4 nsew signal input
rlabel metal2 s 18 0 74 800 6 enc0_b
port 5 nsew signal input
rlabel metal2 s 19338 24752 19394 25552 6 enc1_a
port 6 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 enc1_b
port 7 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 enc2_a
port 8 nsew signal input
rlabel metal3 s 22608 21088 23408 21208 6 enc2_b
port 9 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 pwm0_out
port 10 nsew signal output
rlabel metal2 s 1306 24752 1362 25552 6 pwm1_out
port 11 nsew signal output
rlabel metal2 s 10322 24752 10378 25552 6 pwm2_out
port 12 nsew signal output
rlabel metal3 s 22608 11568 23408 11688 6 reset
port 13 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23408 25552
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1711486
string GDS_FILE /openlane/designs/rgb_mixer/runs/RUN_2025.04.30_22.45.00/results/signoff/rgb_mixer.magic.gds
string GDS_START 312344
<< end >>

