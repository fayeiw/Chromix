* NGSPICE file created from rgb_mixer.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

.subckt rgb_mixer VGND VPWR clk enc0_a enc0_b enc1_a enc1_b enc2_a enc2_b pwm0_out
+ pwm1_out pwm2_out reset
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_501_ _149_ p1.counter\[7\] _165_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_981_ clknet_3_6__leaf_clk _100_ VGND VGND VPWR VPWR e2.value\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_895_ _000_ _001_ VGND VGND VPWR VPWR d0.debounced sky130_fd_sc_hd__dlxtn_1
X_964_ clknet_3_4__leaf_clk _084_ VGND VGND VPWR VPWR d4.state\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_680_ _292_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_878_ net21 _433_ _436_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__o21a_1
X_947_ clknet_3_3__leaf_clk _068_ VGND VGND VPWR VPWR e1.value\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold63 d1.state\[2\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 e0.value\[0\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
Xhold52 p0.counter\[1\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
X_801_ net65 _367_ VGND VGND VPWR VPWR _376_ sky130_fd_sc_hd__and2_1
Xhold41 d3.state\[1\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
X_732_ _331_ _327_ _332_ _308_ VGND VGND VPWR VPWR _333_ sky130_fd_sc_hd__o211ai_2
Xhold74 e1.value\[7\] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
X_663_ net43 _283_ VGND VGND VPWR VPWR _284_ sky130_fd_sc_hd__and2_1
X_594_ _228_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_715_ _317_ _318_ VGND VGND VPWR VPWR _319_ sky130_fd_sc_hd__and2b_1
X_577_ _219_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__clkbuf_1
X_646_ _272_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__clkbuf_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_500_ _149_ p1.counter\[7\] _150_ _164_ VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_629_ _238_ _257_ VGND VGND VPWR VPWR _258_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_980_ clknet_3_6__leaf_clk _099_ VGND VGND VPWR VPWR e2.value\[2\] sky130_fd_sc_hd__dfxtp_1
X_963_ clknet_3_4__leaf_clk _083_ VGND VGND VPWR VPWR d4.state\[3\] sky130_fd_sc_hd__dfxtp_1
X_894_ clknet_3_3__leaf_clk _019_ VGND VGND VPWR VPWR p2.counter\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_877_ _204_ _435_ VGND VGND VPWR VPWR _436_ sky130_fd_sc_hd__nor2_1
X_946_ clknet_3_2__leaf_clk _067_ VGND VGND VPWR VPWR e1.value\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_662_ _201_ VGND VGND VPWR VPWR _283_ sky130_fd_sc_hd__buf_2
Xhold64 d0.state\[5\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 d4.state\[4\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
X_800_ _375_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__clkbuf_1
Xhold53 d6.state\[7\] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 p1.counter\[1\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 d3.state\[7\] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 p1.counter\[5\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
X_731_ e1.value\[4\] _304_ VGND VGND VPWR VPWR _332_ sky130_fd_sc_hd__or2_1
X_593_ net63 _222_ VGND VGND VPWR VPWR _228_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_929_ clknet_3_4__leaf_clk _051_ VGND VGND VPWR VPWR d1.state\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput8 net8 VGND VGND VPWR VPWR pwm0_out sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput10 net10 VGND VGND VPWR VPWR pwm2_out sky130_fd_sc_hd__buf_2
X_645_ _201_ _270_ _271_ VGND VGND VPWR VPWR _272_ sky130_fd_sc_hd__and3_1
X_714_ e1.value\[2\] _303_ VGND VGND VPWR VPWR _318_ sky130_fd_sc_hd__or2_1
X_576_ net69 _212_ VGND VGND VPWR VPWR _219_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_628_ _248_ _246_ _252_ _256_ _247_ VGND VGND VPWR VPWR _257_ sky130_fd_sc_hd__a311o_2
XFILLER_0_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_559_ _204_ _209_ VGND VGND VPWR VPWR _210_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_962_ clknet_3_4__leaf_clk _082_ VGND VGND VPWR VPWR d4.state\[2\] sky130_fd_sc_hd__dfxtp_1
X_893_ clknet_3_3__leaf_clk _018_ VGND VGND VPWR VPWR p2.counter\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_945_ clknet_3_2__leaf_clk _066_ VGND VGND VPWR VPWR e1.value\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_876_ p1.counter\[4\] p1.counter\[3\] _431_ VGND VGND VPWR VPWR _435_ sky130_fd_sc_hd__and3_1
Xhold32 d1.state\[4\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
X_661_ _282_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__clkbuf_1
Xhold76 e0.value\[0\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 d4.state\[7\] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 d5.state\[4\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
X_592_ _227_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__clkbuf_1
Xhold54 d6.state\[5\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 p2.counter\[1\] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 p2.counter\[4\] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlygate4sd3_1
X_730_ e1.value\[4\] _304_ VGND VGND VPWR VPWR _331_ sky130_fd_sc_hd__and2_1
X_928_ clknet_3_4__leaf_clk _050_ VGND VGND VPWR VPWR d1.state\[4\] sky130_fd_sc_hd__dfxtp_1
X_859_ e2.value\[6\] _384_ VGND VGND VPWR VPWR _424_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR pwm1_out sky130_fd_sc_hd__clkbuf_4
X_575_ _218_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__clkbuf_1
X_644_ _236_ _266_ _267_ _269_ VGND VGND VPWR VPWR _271_ sky130_fd_sc_hd__or4_1
X_713_ e1.value\[2\] _303_ VGND VGND VPWR VPWR _317_ sky130_fd_sc_hd__and2_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_627_ e0.value\[3\] _233_ VGND VGND VPWR VPWR _256_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_558_ p2.counter\[6\] p2.counter\[5\] _205_ VGND VGND VPWR VPWR _209_ sky130_fd_sc_hd__and3_1
X_489_ e1.value\[1\] VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_961_ clknet_3_7__leaf_clk _081_ VGND VGND VPWR VPWR d4.state\[1\] sky130_fd_sc_hd__dfxtp_1
X_892_ clknet_3_3__leaf_clk _017_ VGND VGND VPWR VPWR p2.counter\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_944_ clknet_3_3__leaf_clk _065_ VGND VGND VPWR VPWR e1.value\[2\] sky130_fd_sc_hd__dfxtp_1
X_875_ _433_ _434_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold22 _013_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 p1.counter\[4\] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold33 d1.state\[3\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
X_660_ net73 _222_ VGND VGND VPWR VPWR _282_ sky130_fd_sc_hd__and2_1
Xhold55 d5.state\[7\] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlygate4sd3_1
X_591_ net68 _222_ VGND VGND VPWR VPWR _227_ sky130_fd_sc_hd__and2_1
Xhold44 d3.state\[4\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 p1.counter\[3\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_858_ _423_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__clkbuf_1
X_927_ clknet_3_5__leaf_clk _049_ VGND VGND VPWR VPWR d1.state\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_789_ net38 _367_ VGND VGND VPWR VPWR _370_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_712_ e1.value\[1\] _303_ _315_ VGND VGND VPWR VPWR _316_ sky130_fd_sc_hd__o21ba_1
X_574_ net56 _212_ VGND VGND VPWR VPWR _218_ sky130_fd_sc_hd__and2_1
X_643_ _266_ _267_ _269_ _236_ VGND VGND VPWR VPWR _270_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_626_ e0.value\[4\] _233_ VGND VGND VPWR VPWR _255_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_488_ e1.value\[3\] VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__inv_2
X_557_ net29 _205_ _208_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__o21a_1
X_609_ net40 _238_ _240_ VGND VGND VPWR VPWR _241_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_960_ clknet_3_7__leaf_clk _080_ VGND VGND VPWR VPWR d4.state\[0\] sky130_fd_sc_hd__dfxtp_1
X_891_ clknet_3_3__leaf_clk _016_ VGND VGND VPWR VPWR p2.counter\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_943_ clknet_3_3__leaf_clk _064_ VGND VGND VPWR VPWR e1.value\[1\] sky130_fd_sc_hd__dfxtp_1
X_874_ net76 _431_ _202_ VGND VGND VPWR VPWR _434_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold56 d4.state\[5\] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 d6.state\[3\] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 d4.state\[6\] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 d6.state\[4\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold45 p2.counter\[3\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 d0.state\[1\] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
X_590_ _226_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_926_ clknet_3_5__leaf_clk _048_ VGND VGND VPWR VPWR d1.state\[2\] sky130_fd_sc_hd__dfxtp_1
X_788_ _369_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__clkbuf_1
X_857_ _201_ _421_ _422_ VGND VGND VPWR VPWR _423_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_642_ e0.value\[5\] _234_ _257_ _268_ _262_ VGND VGND VPWR VPWR _269_ sky130_fd_sc_hd__a221oi_4
X_711_ _154_ _300_ _313_ _314_ _155_ VGND VGND VPWR VPWR _315_ sky130_fd_sc_hd__o41a_1
X_573_ _217_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_909_ clknet_3_7__leaf_clk _032_ VGND VGND VPWR VPWR d6.state\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_625_ _252_ _253_ _254_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_487_ e1.value\[4\] VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__inv_2
X_556_ _204_ _207_ VGND VGND VPWR VPWR _208_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_608_ _137_ _234_ VGND VGND VPWR VPWR _240_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_539_ net15 _195_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_890_ clknet_3_3__leaf_clk _015_ VGND VGND VPWR VPWR p2.counter\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_942_ clknet_3_0__leaf_clk _063_ VGND VGND VPWR VPWR e1.value\[0\] sky130_fd_sc_hd__dfxtp_1
X_873_ p1.counter\[3\] _431_ VGND VGND VPWR VPWR _433_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold46 d0.state\[6\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 p0.counter\[4\] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 d0.state\[3\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 d4.state\[2\] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 d5.state\[6\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 d3.state\[5\] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
X_925_ clknet_3_5__leaf_clk _047_ VGND VGND VPWR VPWR d1.state\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_787_ _212_ net4 VGND VGND VPWR VPWR _369_ sky130_fd_sc_hd__and2_1
X_856_ _420_ _415_ _416_ _419_ VGND VGND VPWR VPWR _422_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_641_ _255_ _261_ VGND VGND VPWR VPWR _268_ sky130_fd_sc_hd__nor2_1
X_572_ net74 _212_ VGND VGND VPWR VPWR _217_ sky130_fd_sc_hd__and2_1
X_710_ d4.debounced e1.old_a VGND VGND VPWR VPWR _314_ sky130_fd_sc_hd__nor2_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_908_ clknet_3_7__leaf_clk _031_ VGND VGND VPWR VPWR d6.state\[3\] sky130_fd_sc_hd__dfxtp_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_839_ _398_ _396_ _402_ _406_ _397_ VGND VGND VPWR VPWR _407_ sky130_fd_sc_hd__a311o_1
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_624_ _252_ _253_ _195_ VGND VGND VPWR VPWR _254_ sky130_fd_sc_hd__a21oi_1
X_555_ p2.counter\[5\] _205_ VGND VGND VPWR VPWR _207_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_486_ e1.value\[5\] VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_607_ _138_ _236_ _239_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__a21oi_1
X_538_ net7 VGND VGND VPWR VPWR _195_ sky130_fd_sc_hd__buf_4
X_469_ e0.value\[4\] VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_941_ clknet_3_4__leaf_clk _062_ VGND VGND VPWR VPWR e0.old_b sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_872_ _195_ _431_ net26 VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__nor3_1
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold14 d1.state\[6\] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 p0.counter\[2\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 d6.state\[2\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 d5.state\[5\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 d6.state\[6\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 d3.state\[6\] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
X_924_ clknet_3_5__leaf_clk _046_ VGND VGND VPWR VPWR d1.state\[0\] sky130_fd_sc_hd__dfxtp_1
X_786_ _368_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__clkbuf_1
X_855_ _415_ _416_ _419_ _420_ VGND VGND VPWR VPWR _421_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_640_ e0.value\[6\] _234_ VGND VGND VPWR VPWR _267_ sky130_fd_sc_hd__nor2_1
X_571_ _216_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__clkbuf_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_907_ clknet_3_5__leaf_clk _030_ VGND VGND VPWR VPWR d6.state\[2\] sky130_fd_sc_hd__dfxtp_1
X_838_ e2.value\[3\] _383_ VGND VGND VPWR VPWR _406_ sky130_fd_sc_hd__and2_1
X_769_ net17 _356_ _359_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__o21a_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_623_ _247_ _246_ _248_ _238_ VGND VGND VPWR VPWR _253_ sky130_fd_sc_hd__o211a_1
X_554_ net20 _200_ _206_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__o21a_1
X_485_ e1.value\[6\] p1.counter\[6\] VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_468_ e0.value\[5\] VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__inv_2
X_606_ net40 _238_ _196_ VGND VGND VPWR VPWR _239_ sky130_fd_sc_hd__a21o_1
X_537_ _193_ _194_ _010_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_871_ p1.counter\[1\] p1.counter\[0\] net25 VGND VGND VPWR VPWR _432_ sky130_fd_sc_hd__a21oi_1
X_940_ clknet_3_6__leaf_clk _061_ VGND VGND VPWR VPWR d3.state\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold59 d0.state\[7\] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 _351_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 d6.state\[1\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 d4.state\[1\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 p1.counter\[2\] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
X_923_ _004_ _005_ VGND VGND VPWR VPWR d3.debounced sky130_fd_sc_hd__dlxtn_1
X_854_ _384_ _386_ VGND VGND VPWR VPWR _420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_785_ net75 _367_ VGND VGND VPWR VPWR _368_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_570_ net49 _212_ VGND VGND VPWR VPWR _216_ sky130_fd_sc_hd__and2_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_768_ _204_ _358_ VGND VGND VPWR VPWR _359_ sky130_fd_sc_hd__nor2_1
X_906_ clknet_3_5__leaf_clk _029_ VGND VGND VPWR VPWR d6.state\[1\] sky130_fd_sc_hd__dfxtp_1
X_837_ e2.value\[4\] _383_ VGND VGND VPWR VPWR _405_ sky130_fd_sc_hd__xnor2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_699_ _301_ _300_ VGND VGND VPWR VPWR _305_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_622_ _136_ _233_ VGND VGND VPWR VPWR _252_ sky130_fd_sc_hd__xnor2_1
X_553_ _204_ _205_ VGND VGND VPWR VPWR _206_ sky130_fd_sc_hd__nor2_1
X_484_ net84 VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_605_ _237_ VGND VGND VPWR VPWR _238_ sky130_fd_sc_hd__buf_2
X_467_ e0.value\[6\] p0.counter\[6\] VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__and2b_1
X_536_ d6.state\[1\] d6.state\[0\] d6.state\[3\] d6.state\[2\] VGND VGND VPWR VPWR
+ _194_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_519_ e2.value\[7\] _166_ _182_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__a21o_1
XFILLER_0_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_870_ p1.counter\[2\] p1.counter\[1\] p1.counter\[0\] VGND VGND VPWR VPWR _431_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold38 d1.state\[1\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 e1.value\[0\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
Xhold16 _432_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 d5.state\[2\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
X_784_ _201_ VGND VGND VPWR VPWR _367_ sky130_fd_sc_hd__clkbuf_2
X_922_ clknet_3_7__leaf_clk _045_ VGND VGND VPWR VPWR e2.old_b sky130_fd_sc_hd__dfxtp_1
X_853_ _407_ _417_ _418_ VGND VGND VPWR VPWR _419_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_905_ clknet_3_5__leaf_clk _028_ VGND VGND VPWR VPWR d6.state\[0\] sky130_fd_sc_hd__dfxtp_1
X_767_ p0.counter\[6\] p0.counter\[5\] _354_ VGND VGND VPWR VPWR _358_ sky130_fd_sc_hd__and3_1
X_836_ _402_ _403_ _404_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__o21a_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_698_ _303_ VGND VGND VPWR VPWR _304_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_621_ _250_ _251_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__nor2_1
X_483_ _132_ p0.counter\[7\] _148_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__a21oi_1
X_552_ p2.counter\[4\] p2.counter\[3\] _198_ VGND VGND VPWR VPWR _205_ sky130_fd_sc_hd__and3_1
X_819_ _201_ _389_ _390_ VGND VGND VPWR VPWR _391_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_604_ _234_ _235_ VGND VGND VPWR VPWR _237_ sky130_fd_sc_hd__or2_1
X_535_ d6.state\[5\] d6.state\[4\] d6.state\[7\] d6.state\[6\] VGND VGND VPWR VPWR
+ _193_ sky130_fd_sc_hd__or4_1
X_466_ net83 VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_518_ e2.value\[7\] _166_ _167_ _181_ VGND VGND VPWR VPWR _182_ sky130_fd_sc_hd__o22a_1
X_449_ _119_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold39 d0.state\[4\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 d5.state\[1\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 p2.counter\[2\] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd3_1
X_921_ clknet_3_4__leaf_clk _044_ VGND VGND VPWR VPWR e0.old_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_783_ _366_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__clkbuf_1
X_852_ e2.value\[5\] e2.value\[4\] _384_ VGND VGND VPWR VPWR _418_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_904_ clknet_3_5__leaf_clk _027_ VGND VGND VPWR VPWR d0.state\[7\] sky130_fd_sc_hd__dfxtp_1
X_766_ net39 _354_ _357_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__o21a_1
X_697_ _302_ VGND VGND VPWR VPWR _303_ sky130_fd_sc_hd__buf_2
X_835_ _402_ _403_ _259_ VGND VGND VPWR VPWR _404_ sky130_fd_sc_hd__a21oi_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_620_ _238_ _249_ _246_ _196_ VGND VGND VPWR VPWR _251_ sky130_fd_sc_hd__a31o_1
X_551_ _196_ VGND VGND VPWR VPWR _204_ sky130_fd_sc_hd__clkbuf_4
X_482_ _132_ p0.counter\[7\] _133_ _147_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__o22a_1
X_818_ net81 _388_ VGND VGND VPWR VPWR _390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_749_ _343_ _344_ _345_ _347_ _195_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__a311oi_1
X_603_ _234_ _235_ VGND VGND VPWR VPWR _236_ sky130_fd_sc_hd__nor2_2
X_534_ _191_ _192_ _008_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__o21ba_1
X_465_ _131_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_448_ d1.state\[0\] _117_ _118_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_517_ e2.value\[5\] _168_ _178_ _179_ _180_ VGND VGND VPWR VPWR _181_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold29 p0.counter\[5\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 _199_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
X_920_ clknet_3_1__leaf_clk _043_ VGND VGND VPWR VPWR e0.value\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_851_ _405_ _410_ VGND VGND VPWR VPWR _417_ sky130_fd_sc_hd__nor2_1
X_782_ net33 _295_ VGND VGND VPWR VPWR _366_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_903_ clknet_3_5__leaf_clk _026_ VGND VGND VPWR VPWR d0.state\[6\] sky130_fd_sc_hd__dfxtp_1
X_834_ _397_ _396_ _398_ _388_ VGND VGND VPWR VPWR _403_ sky130_fd_sc_hd__o211a_1
X_765_ _204_ _356_ VGND VGND VPWR VPWR _357_ sky130_fd_sc_hd__nor2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_696_ _300_ _301_ VGND VGND VPWR VPWR _302_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_481_ _134_ p0.counter\[5\] _144_ _145_ _146_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__o221a_1
X_550_ _200_ _203_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_817_ e2.value\[0\] _388_ VGND VGND VPWR VPWR _389_ sky130_fd_sc_hd__or2_1
X_679_ net70 _283_ VGND VGND VPWR VPWR _292_ sky130_fd_sc_hd__and2_1
X_748_ _342_ _338_ _346_ _336_ _306_ VGND VGND VPWR VPWR _347_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_602_ _231_ _230_ VGND VGND VPWR VPWR _235_ sky130_fd_sc_hd__and2b_1
X_533_ d5.state\[1\] d5.state\[0\] d5.state\[3\] d5.state\[2\] VGND VGND VPWR VPWR
+ _192_ sky130_fd_sc_hd__or4_1
X_464_ d6.state\[0\] _129_ _130_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_447_ d1.state\[1\] d1.state\[3\] d1.state\[2\] VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_516_ e2.value\[6\] p2.counter\[6\] VGND VGND VPWR VPWR _180_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold19 p2.counter\[5\] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_781_ _365_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__clkbuf_1
X_850_ e2.value\[6\] _384_ VGND VGND VPWR VPWR _416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_979_ clknet_3_3__leaf_clk _098_ VGND VGND VPWR VPWR e2.value\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_902_ clknet_3_5__leaf_clk _025_ VGND VGND VPWR VPWR d0.state\[5\] sky130_fd_sc_hd__dfxtp_1
X_764_ p0.counter\[5\] _354_ VGND VGND VPWR VPWR _356_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_833_ e2.value\[3\] _383_ VGND VGND VPWR VPWR _402_ sky130_fd_sc_hd__xor2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_695_ d4.debounced d3.debounced e1.old_a VGND VGND VPWR VPWR _301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_480_ p0.counter\[6\] e0.value\[6\] VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__or2b_1
X_747_ _344_ _345_ VGND VGND VPWR VPWR _346_ sky130_fd_sc_hd__and2_1
X_816_ _387_ VGND VGND VPWR VPWR _388_ sky130_fd_sc_hd__buf_2
X_678_ _291_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_601_ _233_ VGND VGND VPWR VPWR _234_ sky130_fd_sc_hd__clkbuf_4
X_463_ d6.state\[1\] d6.state\[3\] d6.state\[2\] VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__and3_1
X_532_ d5.state\[5\] d5.state\[4\] d5.state\[7\] d5.state\[6\] VGND VGND VPWR VPWR
+ _191_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_515_ e2.value\[5\] _168_ _169_ e2.value\[4\] VGND VGND VPWR VPWR _179_ sky130_fd_sc_hd__a22o_1
X_446_ d1.state\[5\] d1.state\[4\] d1.state\[7\] d1.state\[6\] VGND VGND VPWR VPWR
+ _117_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 enc0_a VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_780_ net66 _295_ VGND VGND VPWR VPWR _365_ sky130_fd_sc_hd__and2_1
X_978_ clknet_3_6__leaf_clk _097_ VGND VGND VPWR VPWR e2.value\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_901_ clknet_3_5__leaf_clk _024_ VGND VGND VPWR VPWR d0.state\[4\] sky130_fd_sc_hd__dfxtp_1
X_763_ net23 _352_ _355_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__o21a_1
X_694_ d3.debounced d4.debounced e1.old_b VGND VGND VPWR VPWR _300_ sky130_fd_sc_hd__mux2_1
X_832_ _400_ _401_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__nor2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_677_ net61 _283_ VGND VGND VPWR VPWR _291_ sky130_fd_sc_hd__and2_1
X_815_ _384_ _386_ VGND VGND VPWR VPWR _387_ sky130_fd_sc_hd__or2_1
X_746_ _149_ _304_ VGND VGND VPWR VPWR _345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_600_ _232_ VGND VGND VPWR VPWR _233_ sky130_fd_sc_hd__buf_2
X_531_ _189_ _190_ _006_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__o21ba_1
X_462_ d6.state\[5\] d6.state\[4\] d6.state\[7\] d6.state\[6\] VGND VGND VPWR VPWR
+ _129_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_729_ e1.value\[5\] _303_ VGND VGND VPWR VPWR _330_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_514_ e2.value\[4\] _169_ _170_ e2.value\[3\] _177_ VGND VGND VPWR VPWR _178_ sky130_fd_sc_hd__o221a_1
X_445_ _116_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_994_ clknet_3_2__leaf_clk _113_ VGND VGND VPWR VPWR p1.counter\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 enc0_b VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_977_ clknet_3_1__leaf_clk _096_ VGND VGND VPWR VPWR e1.old_b sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_900_ clknet_3_5__leaf_clk _023_ VGND VGND VPWR VPWR d0.state\[3\] sky130_fd_sc_hd__dfxtp_1
X_831_ _388_ _399_ _396_ _196_ VGND VGND VPWR VPWR _401_ sky130_fd_sc_hd__a31o_1
X_762_ _204_ _354_ VGND VGND VPWR VPWR _355_ sky130_fd_sc_hd__nor2_1
X_693_ _299_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__clkbuf_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_814_ _381_ _385_ VGND VGND VPWR VPWR _386_ sky130_fd_sc_hd__and2b_1
X_676_ _290_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__clkbuf_1
X_745_ _149_ _304_ VGND VGND VPWR VPWR _344_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_461_ _128_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__clkbuf_1
X_530_ d4.state\[1\] d4.state\[0\] d4.state\[3\] d4.state\[2\] VGND VGND VPWR VPWR
+ _190_ sky130_fd_sc_hd__or4_1
X_659_ _281_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__clkbuf_1
X_728_ _325_ _328_ _329_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_444_ d0.state\[0\] _114_ _115_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__and3_1
X_513_ _173_ _175_ _176_ VGND VGND VPWR VPWR _177_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_993_ clknet_3_2__leaf_clk _112_ VGND VGND VPWR VPWR p1.counter\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 enc1_a VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_976_ clknet_3_0__leaf_clk _095_ VGND VGND VPWR VPWR d5.state\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_761_ p0.counter\[4\] p0.counter\[3\] _350_ VGND VGND VPWR VPWR _354_ sky130_fd_sc_hd__and3_1
X_830_ _388_ _396_ _399_ VGND VGND VPWR VPWR _400_ sky130_fd_sc_hd__a21oi_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_692_ d1.debounced _295_ VGND VGND VPWR VPWR _299_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_959_ _008_ _009_ VGND VGND VPWR VPWR d5.debounced sky130_fd_sc_hd__dlxtn_1
XFILLER_0_16_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_813_ d5.debounced d6.debounced e2.old_b VGND VGND VPWR VPWR _385_ sky130_fd_sc_hd__mux2_1
X_744_ _342_ _338_ _336_ _306_ VGND VGND VPWR VPWR _343_ sky130_fd_sc_hd__a211o_1
X_675_ net51 _283_ VGND VGND VPWR VPWR _290_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_460_ d5.state\[0\] _126_ _127_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__and3_1
X_727_ _325_ _328_ _259_ VGND VGND VPWR VPWR _329_ sky130_fd_sc_hd__a21oi_1
X_658_ net48 _222_ VGND VGND VPWR VPWR _281_ sky130_fd_sc_hd__and2_1
X_589_ net64 _222_ VGND VGND VPWR VPWR _226_ sky130_fd_sc_hd__and2_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_443_ d0.state\[1\] d0.state\[2\] d0.state\[3\] VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__and3_1
X_512_ e2.value\[3\] _170_ _174_ e2.value\[2\] VGND VGND VPWR VPWR _176_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_992_ clknet_3_2__leaf_clk _111_ VGND VGND VPWR VPWR p1.counter\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput4 enc1_b VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_975_ clknet_3_0__leaf_clk _094_ VGND VGND VPWR VPWR d5.state\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_760_ _352_ _353_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__nor2_1
X_691_ _298_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__clkbuf_1
X_958_ clknet_3_1__leaf_clk _079_ VGND VGND VPWR VPWR p0.counter\[7\] sky130_fd_sc_hd__dfxtp_1
X_889_ clknet_3_3__leaf_clk _014_ VGND VGND VPWR VPWR p2.counter\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_674_ _289_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__clkbuf_1
X_812_ _383_ VGND VGND VPWR VPWR _384_ sky130_fd_sc_hd__buf_2
X_743_ _335_ VGND VGND VPWR VPWR _342_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_657_ _280_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__clkbuf_1
X_726_ _308_ _327_ VGND VGND VPWR VPWR _328_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_588_ _225_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__clkbuf_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_511_ e2.value\[2\] _174_ _171_ e2.value\[1\] VGND VGND VPWR VPWR _175_ sky130_fd_sc_hd__o22a_1
X_442_ d0.state\[4\] d0.state\[5\] d0.state\[6\] d0.state\[7\] VGND VGND VPWR VPWR
+ _114_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_709_ d3.debounced e1.old_a VGND VGND VPWR VPWR _313_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_991_ clknet_3_2__leaf_clk _110_ VGND VGND VPWR VPWR p1.counter\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 enc2_a VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_974_ clknet_3_0__leaf_clk _093_ VGND VGND VPWR VPWR d5.state\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_690_ _202_ net3 VGND VGND VPWR VPWR _298_ sky130_fd_sc_hd__and2_1
X_957_ clknet_3_1__leaf_clk _078_ VGND VGND VPWR VPWR p0.counter\[6\] sky130_fd_sc_hd__dfxtp_1
X_888_ clknet_3_3__leaf_clk net32 VGND VGND VPWR VPWR p2.counter\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_811_ _382_ VGND VGND VPWR VPWR _383_ sky130_fd_sc_hd__clkbuf_2
X_673_ _202_ net2 VGND VGND VPWR VPWR _289_ sky130_fd_sc_hd__and2_1
X_742_ _341_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_587_ net44 _222_ VGND VGND VPWR VPWR _225_ sky130_fd_sc_hd__and2_1
X_656_ d6.debounced _222_ VGND VGND VPWR VPWR _280_ sky130_fd_sc_hd__and2_1
X_725_ _318_ _316_ _322_ _326_ _317_ VGND VGND VPWR VPWR _327_ sky130_fd_sc_hd__a311o_2
XFILLER_0_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_510_ p2.counter\[2\] VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_639_ e0.value\[6\] _234_ VGND VGND VPWR VPWR _266_ sky130_fd_sc_hd__and2_1
X_708_ _311_ _312_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_990_ clknet_3_2__leaf_clk _109_ VGND VGND VPWR VPWR p1.counter\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 enc2_b VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_973_ clknet_3_0__leaf_clk _092_ VGND VGND VPWR VPWR d5.state\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_956_ clknet_3_0__leaf_clk _077_ VGND VGND VPWR VPWR p0.counter\[5\] sky130_fd_sc_hd__dfxtp_1
X_887_ clknet_3_3__leaf_clk _012_ VGND VGND VPWR VPWR p2.counter\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_810_ _379_ _380_ _381_ VGND VGND VPWR VPWR _382_ sky130_fd_sc_hd__and3_1
X_672_ _288_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__clkbuf_1
X_741_ _201_ _339_ _340_ VGND VGND VPWR VPWR _341_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_939_ clknet_3_6__leaf_clk _060_ VGND VGND VPWR VPWR d3.state\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_724_ e1.value\[3\] _303_ VGND VGND VPWR VPWR _326_ sky130_fd_sc_hd__and2_1
X_655_ _279_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__clkbuf_1
X_586_ _224_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_707_ net37 _308_ _310_ _196_ VGND VGND VPWR VPWR _312_ sky130_fd_sc_hd__a31o_1
X_638_ _261_ _264_ _265_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__o21a_1
X_569_ _215_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 reset VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_0_36_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_972_ clknet_3_0__leaf_clk _091_ VGND VGND VPWR VPWR d5.state\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_955_ clknet_3_0__leaf_clk _076_ VGND VGND VPWR VPWR p0.counter\[4\] sky130_fd_sc_hd__dfxtp_1
X_886_ net12 _439_ _441_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_740_ _306_ _335_ _336_ _338_ VGND VGND VPWR VPWR _340_ sky130_fd_sc_hd__or4_1
X_671_ net60 _283_ VGND VGND VPWR VPWR _288_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_869_ net41 net14 _430_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__o21a_1
X_938_ clknet_3_6__leaf_clk _059_ VGND VGND VPWR VPWR d3.state\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_654_ d0.debounced _222_ VGND VGND VPWR VPWR _279_ sky130_fd_sc_hd__and2_1
X_723_ e1.value\[4\] _303_ VGND VGND VPWR VPWR _325_ sky130_fd_sc_hd__xnor2_1
X_585_ net22 _222_ VGND VGND VPWR VPWR _224_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_637_ _261_ _264_ _259_ VGND VGND VPWR VPWR _265_ sky130_fd_sc_hd__a21oi_1
X_706_ net37 _308_ _310_ VGND VGND VPWR VPWR _311_ sky130_fd_sc_hd__a21oi_1
X_568_ net34 _212_ VGND VGND VPWR VPWR _215_ sky130_fd_sc_hd__and2_1
X_499_ _151_ p1.counter\[5\] _161_ _162_ _163_ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_971_ clknet_3_0__leaf_clk _090_ VGND VGND VPWR VPWR d5.state\[2\] sky130_fd_sc_hd__dfxtp_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_954_ clknet_3_1__leaf_clk _075_ VGND VGND VPWR VPWR p0.counter\[3\] sky130_fd_sc_hd__dfxtp_1
X_885_ net12 _439_ _202_ VGND VGND VPWR VPWR _441_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_670_ _287_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__clkbuf_1
X_799_ net45 _367_ VGND VGND VPWR VPWR _375_ sky130_fd_sc_hd__and2_1
X_868_ p1.counter\[1\] p1.counter\[0\] _204_ VGND VGND VPWR VPWR _430_ sky130_fd_sc_hd__a21oi_1
X_937_ clknet_3_6__leaf_clk _058_ VGND VGND VPWR VPWR d3.state\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_653_ _274_ _275_ _276_ _278_ _195_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__a311oi_1
X_722_ _322_ _323_ _324_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__o21a_1
X_584_ _223_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__clkbuf_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_636_ _262_ _257_ _263_ _238_ VGND VGND VPWR VPWR _264_ sky130_fd_sc_hd__o211ai_2
X_567_ _214_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__clkbuf_1
X_705_ _154_ _304_ VGND VGND VPWR VPWR _310_ sky130_fd_sc_hd__xnor2_1
X_498_ p1.counter\[6\] e1.value\[6\] VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__or2b_1
XFILLER_0_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_619_ _238_ _246_ _249_ VGND VGND VPWR VPWR _250_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_970_ clknet_3_0__leaf_clk _089_ VGND VGND VPWR VPWR d5.state\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_953_ clknet_3_0__leaf_clk _074_ VGND VGND VPWR VPWR p0.counter\[2\] sky130_fd_sc_hd__dfxtp_1
X_884_ net16 _437_ _440_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_936_ clknet_3_6__leaf_clk _057_ VGND VGND VPWR VPWR d3.state\[3\] sky130_fd_sc_hd__dfxtp_1
X_798_ _374_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__clkbuf_1
X_867_ net14 _195_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_652_ _273_ _269_ _277_ _267_ _236_ VGND VGND VPWR VPWR _278_ sky130_fd_sc_hd__a2111oi_1
X_583_ net57 _222_ VGND VGND VPWR VPWR _223_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_721_ _322_ _323_ _259_ VGND VGND VPWR VPWR _324_ sky130_fd_sc_hd__a21oi_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_919_ clknet_3_4__leaf_clk _042_ VGND VGND VPWR VPWR e0.value\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 p2.counter\[7\] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_704_ _155_ _306_ _309_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__a21oi_1
X_635_ e0.value\[4\] _234_ VGND VGND VPWR VPWR _263_ sky130_fd_sc_hd__or2_1
X_566_ net72 _212_ VGND VGND VPWR VPWR _214_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_497_ _151_ p1.counter\[5\] p1.counter\[4\] _152_ VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_618_ _247_ _248_ VGND VGND VPWR VPWR _249_ sky130_fd_sc_hd__and2b_1
X_549_ net55 _198_ _202_ VGND VGND VPWR VPWR _203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_952_ clknet_3_0__leaf_clk _073_ VGND VGND VPWR VPWR p0.counter\[1\] sky130_fd_sc_hd__dfxtp_1
X_883_ _204_ _439_ VGND VGND VPWR VPWR _440_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_866_ _429_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__clkbuf_1
X_935_ clknet_3_6__leaf_clk _056_ VGND VGND VPWR VPWR d3.state\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_797_ net46 _367_ VGND VGND VPWR VPWR _374_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_720_ _317_ _316_ _318_ _308_ VGND VGND VPWR VPWR _323_ sky130_fd_sc_hd__o211a_1
X_651_ _275_ _276_ VGND VGND VPWR VPWR _277_ sky130_fd_sc_hd__and2_1
X_582_ _201_ VGND VGND VPWR VPWR _222_ sky130_fd_sc_hd__buf_2
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_918_ clknet_3_1__leaf_clk _041_ VGND VGND VPWR VPWR e0.value\[5\] sky130_fd_sc_hd__dfxtp_1
X_849_ e2.value\[6\] _384_ VGND VGND VPWR VPWR _415_ sky130_fd_sc_hd__and2_1
Xhold2 p1.counter\[7\] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_634_ e0.value\[4\] _234_ VGND VGND VPWR VPWR _262_ sky130_fd_sc_hd__and2_1
X_703_ net37 _308_ _196_ VGND VGND VPWR VPWR _309_ sky130_fd_sc_hd__a21o_1
X_565_ _213_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__clkbuf_1
X_496_ _152_ p1.counter\[4\] p1.counter\[3\] _153_ _160_ VGND VGND VPWR VPWR _161_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_617_ e0.value\[2\] _233_ VGND VGND VPWR VPWR _248_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_479_ _134_ p0.counter\[5\] p0.counter\[4\] _135_ VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__a22o_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_548_ _201_ VGND VGND VPWR VPWR _202_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_951_ clknet_3_0__leaf_clk _072_ VGND VGND VPWR VPWR p0.counter\[0\] sky130_fd_sc_hd__dfxtp_1
X_882_ p1.counter\[6\] p1.counter\[5\] _435_ VGND VGND VPWR VPWR _439_ sky130_fd_sc_hd__and3_1
X_796_ _373_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__clkbuf_1
X_865_ d5.debounced _367_ VGND VGND VPWR VPWR _429_ sky130_fd_sc_hd__and2_1
X_934_ clknet_3_6__leaf_clk _055_ VGND VGND VPWR VPWR d3.state\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_650_ _132_ _234_ VGND VGND VPWR VPWR _276_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_581_ _221_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__clkbuf_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_917_ clknet_3_1__leaf_clk _040_ VGND VGND VPWR VPWR e0.value\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold3 p0.counter\[7\] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlygate4sd3_1
X_779_ _364_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__clkbuf_1
X_848_ _410_ _413_ _414_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__o21a_1
X_633_ e0.value\[5\] _233_ VGND VGND VPWR VPWR _261_ sky130_fd_sc_hd__xnor2_1
X_702_ _307_ VGND VGND VPWR VPWR _308_ sky130_fd_sc_hd__buf_2
X_564_ net77 _212_ VGND VGND VPWR VPWR _213_ sky130_fd_sc_hd__and2_1
X_495_ _156_ _158_ _159_ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_616_ e0.value\[2\] _233_ VGND VGND VPWR VPWR _247_ sky130_fd_sc_hd__and2_1
X_547_ net7 VGND VGND VPWR VPWR _201_ sky130_fd_sc_hd__inv_2
X_478_ _135_ p0.counter\[4\] p0.counter\[3\] _136_ _143_ VGND VGND VPWR VPWR _144_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_950_ clknet_3_3__leaf_clk _071_ VGND VGND VPWR VPWR e1.old_a sky130_fd_sc_hd__dfxtp_1
X_881_ net30 _435_ _438_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_933_ clknet_3_7__leaf_clk _054_ VGND VGND VPWR VPWR d3.state\[0\] sky130_fd_sc_hd__dfxtp_1
X_795_ net53 _367_ VGND VGND VPWR VPWR _373_ sky130_fd_sc_hd__and2_1
X_864_ _195_ _427_ _428_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__nor3b_1
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_580_ net47 _212_ VGND VGND VPWR VPWR _221_ sky130_fd_sc_hd__and2_1
X_916_ clknet_3_1__leaf_clk _039_ VGND VGND VPWR VPWR e0.value\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold4 p1.counter\[0\] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_778_ net52 _295_ VGND VGND VPWR VPWR _364_ sky130_fd_sc_hd__and2_1
X_847_ _410_ _413_ _259_ VGND VGND VPWR VPWR _414_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_632_ _255_ _258_ _260_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__o21a_1
X_563_ _201_ VGND VGND VPWR VPWR _212_ sky130_fd_sc_hd__buf_2
X_701_ _304_ _305_ VGND VGND VPWR VPWR _307_ sky130_fd_sc_hd__or2_1
X_494_ _153_ p1.counter\[3\] p1.counter\[2\] _157_ VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_615_ e0.value\[1\] _233_ _245_ VGND VGND VPWR VPWR _246_ sky130_fd_sc_hd__o21ba_1
X_546_ p2.counter\[3\] _198_ VGND VGND VPWR VPWR _200_ sky130_fd_sc_hd__and2_1
X_477_ _139_ _141_ _142_ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_529_ d4.state\[5\] d4.state\[4\] d4.state\[7\] d4.state\[6\] VGND VGND VPWR VPWR
+ _189_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_880_ _204_ _437_ VGND VGND VPWR VPWR _438_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_932_ _006_ _007_ VGND VGND VPWR VPWR d4.debounced sky130_fd_sc_hd__dlxtn_1
X_863_ _388_ _424_ _425_ _426_ VGND VGND VPWR VPWR _428_ sky130_fd_sc_hd__a31o_1
X_794_ _372_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_915_ clknet_3_1__leaf_clk _038_ VGND VGND VPWR VPWR e0.value\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold5 p2.counter\[0\] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlygate4sd3_1
X_846_ _411_ _407_ _412_ _388_ VGND VGND VPWR VPWR _413_ sky130_fd_sc_hd__o211ai_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_777_ _363_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_700_ _304_ _305_ VGND VGND VPWR VPWR _306_ sky130_fd_sc_hd__nor2_2
X_631_ _255_ _258_ _259_ VGND VGND VPWR VPWR _260_ sky130_fd_sc_hd__a21oi_1
X_493_ _157_ p1.counter\[2\] p1.counter\[1\] _154_ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__o22a_1
X_562_ net11 _209_ _211_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_829_ _397_ _398_ VGND VGND VPWR VPWR _399_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_476_ _136_ p0.counter\[3\] p0.counter\[2\] _140_ VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__a22o_1
X_614_ _137_ _230_ _243_ _244_ _138_ VGND VGND VPWR VPWR _245_ sky130_fd_sc_hd__o41a_1
X_545_ _195_ _198_ net28 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__nor3_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_459_ d5.state\[1\] d5.state\[3\] d5.state\[2\] VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__and3_1
X_528_ _187_ _188_ _004_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_23_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_931_ clknet_3_4__leaf_clk _053_ VGND VGND VPWR VPWR d1.state\[7\] sky130_fd_sc_hd__dfxtp_1
X_862_ _388_ _424_ _425_ _426_ VGND VGND VPWR VPWR _427_ sky130_fd_sc_hd__and4_1
X_793_ net82 _367_ VGND VGND VPWR VPWR _372_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_914_ clknet_3_4__leaf_clk _037_ VGND VGND VPWR VPWR e0.value\[1\] sky130_fd_sc_hd__dfxtp_1
X_776_ net50 _295_ VGND VGND VPWR VPWR _363_ sky130_fd_sc_hd__and2_1
X_845_ e2.value\[4\] _384_ VGND VGND VPWR VPWR _412_ sky130_fd_sc_hd__or2_1
Xhold6 p1.counter\[6\] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_630_ _196_ VGND VGND VPWR VPWR _259_ sky130_fd_sc_hd__clkbuf_4
X_492_ e1.value\[2\] VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__inv_2
X_561_ net11 _209_ _202_ VGND VGND VPWR VPWR _211_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_759_ net80 _350_ _202_ VGND VGND VPWR VPWR _353_ sky130_fd_sc_hd__o21ai_1
X_828_ e2.value\[2\] _383_ VGND VGND VPWR VPWR _398_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_613_ d1.debounced e0.old_a VGND VGND VPWR VPWR _244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_475_ _140_ p0.counter\[2\] p0.counter\[1\] _137_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__o22a_1
X_544_ p2.counter\[1\] p2.counter\[0\] net27 VGND VGND VPWR VPWR _199_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_527_ d3.state\[1\] d3.state\[0\] d3.state\[3\] d3.state\[2\] VGND VGND VPWR VPWR
+ _188_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_458_ d5.state\[5\] d5.state\[4\] d5.state\[7\] d5.state\[6\] VGND VGND VPWR VPWR
+ _126_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_930_ clknet_3_5__leaf_clk _052_ VGND VGND VPWR VPWR d1.state\[6\] sky130_fd_sc_hd__dfxtp_1
X_792_ _371_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__clkbuf_1
X_861_ e2.value\[7\] _384_ VGND VGND VPWR VPWR _426_ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_913_ clknet_3_4__leaf_clk _036_ VGND VGND VPWR VPWR e0.value\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold7 p0.counter\[6\] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlygate4sd3_1
X_775_ _362_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__clkbuf_1
X_844_ e2.value\[4\] _384_ VGND VGND VPWR VPWR _411_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_560_ net19 _207_ _210_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__o21a_1
X_491_ _154_ p1.counter\[1\] p1.counter\[0\] _155_ VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_758_ p0.counter\[3\] _350_ VGND VGND VPWR VPWR _352_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_689_ _297_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__clkbuf_1
X_827_ e2.value\[2\] _383_ VGND VGND VPWR VPWR _397_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_612_ d0.debounced e0.old_a VGND VGND VPWR VPWR _243_ sky130_fd_sc_hd__and2b_1
X_543_ p2.counter\[2\] p2.counter\[1\] p2.counter\[0\] VGND VGND VPWR VPWR _198_ sky130_fd_sc_hd__and3_1
X_474_ e0.value\[2\] VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_526_ d3.state\[5\] d3.state\[4\] d3.state\[7\] d3.state\[6\] VGND VGND VPWR VPWR
+ _187_ sky130_fd_sc_hd__or4_1
X_457_ _125_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_509_ e2.value\[1\] _171_ _172_ e2.value\[0\] VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__a22o_1
X_791_ net59 _367_ VGND VGND VPWR VPWR _371_ sky130_fd_sc_hd__and2_1
X_860_ _407_ _417_ _418_ _415_ VGND VGND VPWR VPWR _425_ sky130_fd_sc_hd__a211o_1
X_989_ clknet_3_2__leaf_clk _108_ VGND VGND VPWR VPWR p1.counter\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_912_ clknet_3_7__leaf_clk _035_ VGND VGND VPWR VPWR d6.state\[7\] sky130_fd_sc_hd__dfxtp_1
X_843_ e2.value\[5\] _384_ VGND VGND VPWR VPWR _410_ sky130_fd_sc_hd__xnor2_1
Xhold8 p0.counter\[0\] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlygate4sd3_1
X_774_ net78 _295_ VGND VGND VPWR VPWR _362_ sky130_fd_sc_hd__and2_1
X_490_ net37 VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_826_ e2.value\[0\] _392_ _393_ VGND VGND VPWR VPWR _396_ sky130_fd_sc_hd__o21a_1
X_757_ _195_ _350_ net36 VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__nor3_1
XFILLER_0_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_688_ net85 _295_ VGND VGND VPWR VPWR _297_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_473_ _137_ p0.counter\[1\] p0.counter\[0\] _138_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__a211o_1
X_611_ _241_ _242_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__nor2_1
X_542_ _171_ _172_ _197_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_809_ d6.debounced d5.debounced e2.old_a VGND VGND VPWR VPWR _381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_525_ _185_ _186_ _002_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__o21ba_1
X_456_ d4.state\[0\] _123_ _124_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_508_ net15 VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_790_ _370_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__clkbuf_1
X_988_ clknet_3_2__leaf_clk _107_ VGND VGND VPWR VPWR p1.counter\[1\] sky130_fd_sc_hd__dfxtp_1
X_911_ clknet_3_7__leaf_clk _034_ VGND VGND VPWR VPWR d6.state\[6\] sky130_fd_sc_hd__dfxtp_1
X_842_ _405_ _408_ _409_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__o21a_1
Xhold9 p2.counter\[6\] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlygate4sd3_1
X_773_ _361_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_756_ p0.counter\[0\] p0.counter\[1\] net35 VGND VGND VPWR VPWR _351_ sky130_fd_sc_hd__a21oi_1
X_825_ _390_ _394_ _395_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__o21a_1
X_687_ _296_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_610_ net86 _238_ _240_ _196_ VGND VGND VPWR VPWR _242_ sky130_fd_sc_hd__a31o_1
X_472_ net40 VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__inv_2
X_541_ net31 p2.counter\[0\] _196_ VGND VGND VPWR VPWR _197_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_808_ d6.debounced e2.old_b VGND VGND VPWR VPWR _380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_739_ _335_ _336_ _338_ _306_ VGND VGND VPWR VPWR _339_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_524_ d1.state\[1\] d1.state\[0\] d1.state\[3\] d1.state\[2\] VGND VGND VPWR VPWR
+ _186_ sky130_fd_sc_hd__or4_1
X_455_ d4.state\[1\] d4.state\[3\] d4.state\[2\] VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_507_ net31 VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_987_ clknet_3_0__leaf_clk _106_ VGND VGND VPWR VPWR p1.counter\[0\] sky130_fd_sc_hd__dfxtp_1
X_772_ net58 _295_ VGND VGND VPWR VPWR _361_ sky130_fd_sc_hd__and2_1
X_910_ clknet_3_7__leaf_clk _033_ VGND VGND VPWR VPWR d6.state\[5\] sky130_fd_sc_hd__dfxtp_1
X_841_ _405_ _408_ _259_ VGND VGND VPWR VPWR _409_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_755_ p0.counter\[0\] p0.counter\[2\] p0.counter\[1\] VGND VGND VPWR VPWR _350_ sky130_fd_sc_hd__and3_1
X_824_ _390_ _394_ _259_ VGND VGND VPWR VPWR _395_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_686_ net79 _295_ VGND VGND VPWR VPWR _296_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_540_ net7 VGND VGND VPWR VPWR _196_ sky130_fd_sc_hd__clkbuf_4
X_471_ e0.value\[1\] VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__inv_2
X_669_ net24 _283_ VGND VGND VPWR VPWR _287_ sky130_fd_sc_hd__and2_1
X_807_ e2.old_b d5.debounced VGND VGND VPWR VPWR _379_ sky130_fd_sc_hd__or2b_1
X_738_ e1.value\[5\] _304_ _327_ _337_ _331_ VGND VGND VPWR VPWR _338_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_523_ d1.state\[5\] d1.state\[4\] d1.state\[7\] d1.state\[6\] VGND VGND VPWR VPWR
+ _185_ sky130_fd_sc_hd__or4_1
X_454_ d4.state\[5\] d4.state\[4\] d4.state\[7\] d4.state\[6\] VGND VGND VPWR VPWR
+ _123_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_506_ p2.counter\[3\] VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_986_ clknet_3_3__leaf_clk _105_ VGND VGND VPWR VPWR e2.old_a sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_771_ net13 _358_ _360_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__a21oi_1
X_840_ _388_ _407_ VGND VGND VPWR VPWR _408_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_969_ clknet_3_1__leaf_clk _088_ VGND VGND VPWR VPWR d5.state\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_823_ _392_ _393_ VGND VGND VPWR VPWR _394_ sky130_fd_sc_hd__or2b_1
X_754_ net18 net62 _349_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__o21a_1
X_685_ _201_ VGND VGND VPWR VPWR _295_ sky130_fd_sc_hd__buf_2
XFILLER_0_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_470_ e0.value\[3\] VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__inv_2
X_806_ _378_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__clkbuf_1
X_599_ _230_ _231_ VGND VGND VPWR VPWR _232_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_668_ _286_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__clkbuf_1
X_737_ _325_ _330_ VGND VGND VPWR VPWR _337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_522_ _183_ _184_ _000_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__o21ba_1
X_453_ _122_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_505_ p2.counter\[4\] VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_985_ clknet_3_6__leaf_clk _104_ VGND VGND VPWR VPWR e2.value\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_770_ net13 _358_ _202_ VGND VGND VPWR VPWR _360_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_968_ _010_ _011_ VGND VGND VPWR VPWR d6.debounced sky130_fd_sc_hd__dlxtn_1
XFILLER_0_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_899_ clknet_3_4__leaf_clk _022_ VGND VGND VPWR VPWR d0.state\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_822_ _379_ _380_ _381_ e2.value\[1\] VGND VGND VPWR VPWR _393_ sky130_fd_sc_hd__a31o_1
X_753_ p0.counter\[0\] p0.counter\[1\] _259_ VGND VGND VPWR VPWR _349_ sky130_fd_sc_hd__a21oi_1
X_684_ _294_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__clkbuf_1
Xhold70 p0.counter\[3\] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
X_805_ d4.debounced _367_ VGND VGND VPWR VPWR _378_ sky130_fd_sc_hd__and2_1
X_736_ e1.value\[6\] _304_ VGND VGND VPWR VPWR _336_ sky130_fd_sc_hd__nor2_1
X_598_ d1.debounced d0.debounced e0.old_a VGND VGND VPWR VPWR _231_ sky130_fd_sc_hd__mux2_1
X_667_ net71 _283_ VGND VGND VPWR VPWR _286_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_521_ d0.state\[0\] d0.state\[1\] d0.state\[2\] d0.state\[3\] VGND VGND VPWR VPWR
+ _184_ sky130_fd_sc_hd__or4_1
X_452_ d3.state\[0\] _120_ _121_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_719_ _153_ _303_ VGND VGND VPWR VPWR _322_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_504_ p2.counter\[5\] VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_984_ clknet_3_6__leaf_clk _103_ VGND VGND VPWR VPWR e2.value\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_898_ clknet_3_4__leaf_clk _021_ VGND VGND VPWR VPWR d0.state\[1\] sky130_fd_sc_hd__dfxtp_1
X_967_ clknet_3_4__leaf_clk _087_ VGND VGND VPWR VPWR d4.state\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_752_ net18 _195_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__nor2_1
X_821_ _385_ _381_ e2.value\[1\] VGND VGND VPWR VPWR _392_ sky130_fd_sc_hd__and3b_1
X_683_ net67 _283_ VGND VGND VPWR VPWR _294_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_804_ _377_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__clkbuf_1
Xhold71 e2.value\[0\] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold60 d3.state\[3\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
X_735_ e1.value\[6\] _304_ VGND VGND VPWR VPWR _335_ sky130_fd_sc_hd__and2_1
X_666_ _285_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__clkbuf_1
X_597_ d0.debounced d1.debounced e0.old_b VGND VGND VPWR VPWR _230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_520_ d0.state\[4\] d0.state\[5\] d0.state\[6\] d0.state\[7\] VGND VGND VPWR VPWR
+ _183_ sky130_fd_sc_hd__or4_1
X_451_ d3.state\[1\] d3.state\[3\] d3.state\[2\] VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_649_ _132_ _234_ VGND VGND VPWR VPWR _275_ sky130_fd_sc_hd__or2_1
X_718_ _320_ _321_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_503_ p2.counter\[6\] e2.value\[6\] VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_983_ clknet_3_6__leaf_clk _102_ VGND VGND VPWR VPWR e2.value\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_897_ clknet_3_4__leaf_clk _020_ VGND VGND VPWR VPWR d0.state\[0\] sky130_fd_sc_hd__dfxtp_1
X_966_ clknet_3_1__leaf_clk _086_ VGND VGND VPWR VPWR d4.state\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_751_ _348_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__clkbuf_1
X_820_ _391_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__clkbuf_1
X_682_ _293_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__clkbuf_1
X_949_ clknet_3_2__leaf_clk _070_ VGND VGND VPWR VPWR e1.value\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_665_ net42 _283_ VGND VGND VPWR VPWR _285_ sky130_fd_sc_hd__and2_1
Xhold50 d1.state\[7\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 d1.state\[5\] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
X_803_ _212_ net5 VGND VGND VPWR VPWR _377_ sky130_fd_sc_hd__and2_1
Xhold72 d5.state\[3\] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
X_734_ _330_ _333_ _334_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__o21a_1
X_596_ _229_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_450_ d3.state\[5\] d3.state\[4\] d3.state\[7\] d3.state\[6\] VGND VGND VPWR VPWR
+ _120_ sky130_fd_sc_hd__and4_1
X_648_ _273_ _269_ _267_ _236_ VGND VGND VPWR VPWR _274_ sky130_fd_sc_hd__a211o_1
X_717_ _308_ _319_ _316_ _196_ VGND VGND VPWR VPWR _321_ sky130_fd_sc_hd__a31o_1
X_579_ _220_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__clkbuf_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_502_ p2.counter\[7\] VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_982_ clknet_3_6__leaf_clk _101_ VGND VGND VPWR VPWR e2.value\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_965_ clknet_3_4__leaf_clk _085_ VGND VGND VPWR VPWR d4.state\[5\] sky130_fd_sc_hd__dfxtp_1
X_896_ _002_ _003_ VGND VGND VPWR VPWR d1.debounced sky130_fd_sc_hd__dlxtn_1
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_750_ d3.debounced _295_ VGND VGND VPWR VPWR _348_ sky130_fd_sc_hd__and2_1
X_681_ net54 _283_ VGND VGND VPWR VPWR _293_ sky130_fd_sc_hd__and2_1
X_948_ clknet_3_3__leaf_clk _069_ VGND VGND VPWR VPWR e1.value\[6\] sky130_fd_sc_hd__dfxtp_1
X_879_ p1.counter\[5\] _435_ VGND VGND VPWR VPWR _437_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_802_ _376_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__clkbuf_1
Xhold40 d4.state\[3\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_664_ _284_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__clkbuf_1
Xhold62 d0.state\[2\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 e0.value\[7\] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 d3.state\[2\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
X_733_ _330_ _333_ _259_ VGND VGND VPWR VPWR _334_ sky130_fd_sc_hd__a21oi_1
X_595_ _202_ net6 VGND VGND VPWR VPWR _229_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_716_ _308_ _316_ _319_ VGND VGND VPWR VPWR _320_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_647_ _266_ VGND VGND VPWR VPWR _273_ sky130_fd_sc_hd__inv_2
X_578_ _202_ net1 VGND VGND VPWR VPWR _220_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

