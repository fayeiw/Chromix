magic
tech sky130A
magscale 1 2
timestamp 1746053288
<< checkpaint >>
rect -1260 7244 24668 26812
rect -2866 -1260 24668 7244
<< viali >>
rect 1501 22729 1535 22763
rect 10701 22729 10735 22763
rect 1777 22593 1811 22627
rect 10885 22593 10919 22627
rect 13277 22593 13311 22627
rect 13461 22593 13495 22627
rect 13645 22593 13679 22627
rect 13737 22593 13771 22627
rect 16773 22593 16807 22627
rect 19625 22593 19659 22627
rect 16957 22389 16991 22423
rect 19441 22389 19475 22423
rect 7481 22185 7515 22219
rect 7389 22117 7423 22151
rect 13553 22117 13587 22151
rect 5181 22049 5215 22083
rect 7481 22049 7515 22083
rect 13277 22049 13311 22083
rect 3249 21981 3283 22015
rect 4353 21981 4387 22015
rect 7297 21981 7331 22015
rect 7757 21981 7791 22015
rect 8309 21981 8343 22015
rect 9965 21981 9999 22015
rect 11989 21981 12023 22015
rect 12449 21981 12483 22015
rect 13093 21981 13127 22015
rect 15485 21981 15519 22015
rect 17877 21981 17911 22015
rect 2973 21913 3007 21947
rect 5448 21913 5482 21947
rect 7665 21913 7699 21947
rect 10232 21913 10266 21947
rect 12173 21913 12207 21947
rect 12357 21913 12391 21947
rect 12541 21913 12575 21947
rect 15218 21913 15252 21947
rect 17610 21913 17644 21947
rect 3071 21845 3105 21879
rect 3157 21845 3191 21879
rect 3801 21845 3835 21879
rect 6561 21845 6595 21879
rect 7849 21845 7883 21879
rect 8493 21845 8527 21879
rect 11345 21845 11379 21879
rect 11437 21845 11471 21879
rect 12271 21845 12305 21879
rect 13737 21845 13771 21879
rect 14105 21845 14139 21879
rect 16497 21845 16531 21879
rect 5733 21641 5767 21675
rect 6009 21641 6043 21675
rect 6929 21641 6963 21675
rect 10425 21641 10459 21675
rect 13093 21641 13127 21675
rect 13185 21641 13219 21675
rect 14289 21641 14323 21675
rect 17141 21641 17175 21675
rect 17391 21641 17425 21675
rect 2964 21573 2998 21607
rect 5181 21573 5215 21607
rect 6101 21573 6135 21607
rect 9146 21573 9180 21607
rect 11980 21573 12014 21607
rect 15209 21573 15243 21607
rect 17601 21573 17635 21607
rect 2329 21505 2363 21539
rect 2513 21505 2547 21539
rect 2605 21505 2639 21539
rect 5365 21505 5399 21539
rect 5549 21505 5583 21539
rect 5733 21505 5767 21539
rect 6193 21505 6227 21539
rect 6561 21505 6595 21539
rect 6837 21505 6871 21539
rect 7665 21505 7699 21539
rect 10609 21505 10643 21539
rect 10885 21505 10919 21539
rect 10977 21505 11011 21539
rect 11161 21505 11195 21539
rect 13369 21505 13403 21539
rect 13461 21505 13495 21539
rect 13737 21505 13771 21539
rect 14565 21505 14599 21539
rect 15025 21505 15059 21539
rect 15853 21505 15887 21539
rect 16037 21505 16071 21539
rect 16129 21505 16163 21539
rect 16497 21505 16531 21539
rect 16681 21505 16715 21539
rect 16957 21505 16991 21539
rect 21649 21505 21683 21539
rect 2697 21437 2731 21471
rect 6653 21437 6687 21471
rect 9413 21437 9447 21471
rect 11069 21437 11103 21471
rect 11713 21437 11747 21471
rect 13921 21437 13955 21471
rect 14013 21437 14047 21471
rect 14105 21437 14139 21471
rect 14657 21437 14691 21471
rect 16313 21437 16347 21471
rect 16773 21437 16807 21471
rect 2329 21369 2363 21403
rect 4077 21369 4111 21403
rect 8033 21369 8067 21403
rect 13645 21369 13679 21403
rect 16037 21369 16071 21403
rect 16221 21369 16255 21403
rect 5825 21301 5859 21335
rect 6377 21301 6411 21335
rect 6745 21301 6779 21335
rect 7113 21301 7147 21335
rect 10793 21301 10827 21335
rect 14933 21301 14967 21335
rect 15393 21301 15427 21335
rect 16313 21301 16347 21335
rect 16773 21301 16807 21335
rect 17233 21301 17267 21335
rect 17417 21301 17451 21335
rect 21465 21301 21499 21335
rect 3341 21097 3375 21131
rect 3433 21097 3467 21131
rect 3801 21097 3835 21131
rect 4261 21097 4295 21131
rect 6377 21097 6411 21131
rect 7021 21097 7055 21131
rect 7757 21097 7791 21131
rect 8309 21097 8343 21131
rect 8493 21097 8527 21131
rect 9689 21097 9723 21131
rect 11989 21097 12023 21131
rect 12173 21097 12207 21131
rect 13001 21097 13035 21131
rect 13369 21097 13403 21131
rect 14749 21097 14783 21131
rect 15393 21097 15427 21131
rect 17049 21097 17083 21131
rect 5825 21029 5859 21063
rect 7113 21029 7147 21063
rect 11161 21029 11195 21063
rect 3249 20961 3283 20995
rect 6009 20961 6043 20995
rect 6653 20961 6687 20995
rect 7849 20961 7883 20995
rect 11897 20961 11931 20995
rect 15669 20961 15703 20995
rect 15761 20961 15795 20995
rect 16681 20961 16715 20995
rect 3525 20893 3559 20927
rect 3985 20893 4019 20927
rect 4077 20893 4111 20927
rect 4353 20893 4387 20927
rect 5733 20893 5767 20927
rect 5917 20893 5951 20927
rect 6193 20893 6227 20927
rect 6837 20893 6871 20927
rect 7311 20871 7345 20905
rect 7462 20893 7496 20927
rect 7573 20893 7607 20927
rect 7665 20893 7699 20927
rect 8033 20893 8067 20927
rect 9505 20893 9539 20927
rect 9689 20893 9723 20927
rect 9781 20893 9815 20927
rect 12725 20893 12759 20927
rect 13277 20893 13311 20927
rect 14933 20893 14967 20927
rect 15025 20893 15059 20927
rect 15117 20893 15151 20927
rect 15577 20893 15611 20927
rect 15853 20893 15887 20927
rect 16865 20893 16899 20927
rect 7757 20825 7791 20859
rect 8677 20825 8711 20859
rect 10048 20825 10082 20859
rect 12141 20825 12175 20859
rect 12357 20825 12391 20859
rect 15301 20825 15335 20859
rect 8217 20757 8251 20791
rect 8467 20757 8501 20791
rect 11253 20757 11287 20791
rect 13185 20757 13219 20791
rect 3893 20553 3927 20587
rect 6561 20553 6595 20587
rect 6837 20553 6871 20587
rect 10241 20553 10275 20587
rect 10793 20553 10827 20587
rect 11989 20553 12023 20587
rect 15301 20553 15335 20587
rect 15853 20553 15887 20587
rect 9045 20485 9079 20519
rect 6653 20417 6687 20451
rect 6745 20417 6779 20451
rect 6929 20417 6963 20451
rect 10425 20417 10459 20451
rect 10977 20417 11011 20451
rect 12173 20417 12207 20451
rect 12265 20417 12299 20451
rect 12449 20417 12483 20451
rect 15209 20417 15243 20451
rect 15393 20417 15427 20451
rect 15761 20417 15795 20451
rect 16037 20417 16071 20451
rect 16129 20417 16163 20451
rect 16313 20417 16347 20451
rect 16405 20417 16439 20451
rect 16681 20417 16715 20451
rect 16865 20417 16899 20451
rect 16957 20417 16991 20451
rect 20361 20417 20395 20451
rect 3433 20349 3467 20383
rect 10701 20349 10735 20383
rect 11161 20349 11195 20383
rect 11989 20349 12023 20383
rect 20177 20349 20211 20383
rect 3801 20281 3835 20315
rect 16681 20281 16715 20315
rect 9137 20213 9171 20247
rect 10609 20213 10643 20247
rect 12541 20213 12575 20247
rect 15577 20213 15611 20247
rect 20545 20213 20579 20247
rect 4721 20009 4755 20043
rect 13737 20009 13771 20043
rect 15761 20009 15795 20043
rect 16405 20009 16439 20043
rect 16773 20009 16807 20043
rect 13369 19873 13403 19907
rect 16865 19873 16899 19907
rect 17693 19873 17727 19907
rect 19625 19873 19659 19907
rect 2881 19805 2915 19839
rect 3065 19805 3099 19839
rect 3157 19805 3191 19839
rect 3341 19805 3375 19839
rect 4353 19805 4387 19839
rect 4997 19805 5031 19839
rect 13001 19805 13035 19839
rect 13185 19805 13219 19839
rect 13277 19805 13311 19839
rect 13553 19805 13587 19839
rect 15577 19805 15611 19839
rect 16589 19805 16623 19839
rect 17601 19805 17635 19839
rect 19441 19805 19475 19839
rect 20453 19805 20487 19839
rect 15393 19737 15427 19771
rect 2973 19669 3007 19703
rect 3249 19669 3283 19703
rect 3801 19669 3835 19703
rect 4537 19669 4571 19703
rect 17969 19669 18003 19703
rect 19257 19669 19291 19703
rect 20269 19669 20303 19703
rect 2789 19465 2823 19499
rect 3433 19465 3467 19499
rect 13461 19465 13495 19499
rect 17693 19465 17727 19499
rect 3601 19397 3635 19431
rect 3801 19397 3835 19431
rect 6009 19397 6043 19431
rect 12725 19397 12759 19431
rect 13093 19397 13127 19431
rect 13185 19397 13219 19431
rect 1409 19329 1443 19363
rect 1676 19329 1710 19363
rect 2881 19329 2915 19363
rect 3065 19329 3099 19363
rect 3341 19329 3375 19363
rect 5917 19329 5951 19363
rect 6193 19329 6227 19363
rect 6561 19329 6595 19363
rect 6837 19329 6871 19363
rect 7021 19329 7055 19363
rect 7297 19329 7331 19363
rect 7481 19329 7515 19363
rect 8125 19329 8159 19363
rect 10333 19329 10367 19363
rect 10517 19329 10551 19363
rect 11069 19329 11103 19363
rect 11897 19329 11931 19363
rect 12633 19329 12667 19363
rect 12909 19329 12943 19363
rect 13277 19329 13311 19363
rect 16313 19329 16347 19363
rect 16497 19329 16531 19363
rect 16669 19351 16703 19385
rect 16773 19329 16807 19363
rect 17417 19329 17451 19363
rect 17601 19329 17635 19363
rect 18806 19329 18840 19363
rect 19073 19329 19107 19363
rect 19165 19329 19199 19363
rect 6377 19261 6411 19295
rect 8401 19261 8435 19295
rect 11253 19261 11287 19295
rect 12449 19261 12483 19295
rect 16129 19261 16163 19295
rect 16957 19261 16991 19295
rect 17049 19261 17083 19295
rect 17233 19193 17267 19227
rect 3249 19125 3283 19159
rect 3617 19125 3651 19159
rect 6193 19125 6227 19159
rect 6745 19125 6779 19159
rect 7205 19125 7239 19159
rect 7481 19125 7515 19159
rect 7941 19125 7975 19159
rect 8309 19125 8343 19159
rect 10517 19125 10551 19159
rect 10885 19125 10919 19159
rect 17141 19125 17175 19159
rect 19349 19125 19383 19159
rect 3801 18921 3835 18955
rect 9229 18921 9263 18955
rect 10333 18921 10367 18955
rect 11897 18921 11931 18955
rect 12173 18921 12207 18955
rect 16037 18921 16071 18955
rect 16865 18921 16899 18955
rect 17509 18921 17543 18955
rect 17877 18921 17911 18955
rect 7297 18853 7331 18887
rect 17969 18853 18003 18887
rect 2237 18785 2271 18819
rect 4721 18785 4755 18819
rect 4905 18785 4939 18819
rect 10517 18785 10551 18819
rect 15485 18785 15519 18819
rect 3985 18717 4019 18751
rect 4169 18717 4203 18751
rect 4261 18717 4295 18751
rect 4353 18717 4387 18751
rect 4537 18717 4571 18751
rect 4813 18717 4847 18751
rect 6745 18717 6779 18751
rect 7113 18717 7147 18751
rect 7389 18717 7423 18751
rect 7656 18717 7690 18751
rect 8953 18717 8987 18751
rect 9045 18717 9079 18751
rect 10149 18717 10183 18751
rect 10425 18717 10459 18751
rect 13921 18717 13955 18751
rect 15393 18717 15427 18751
rect 15853 18717 15887 18751
rect 16681 18717 16715 18751
rect 16865 18717 16899 18751
rect 17417 18717 17451 18751
rect 17693 18717 17727 18751
rect 18153 18717 18187 18751
rect 18245 18717 18279 18751
rect 20637 18717 20671 18751
rect 12127 18683 12161 18717
rect 2504 18649 2538 18683
rect 5172 18649 5206 18683
rect 6469 18649 6503 18683
rect 7205 18649 7239 18683
rect 9229 18649 9263 18683
rect 10784 18649 10818 18683
rect 12357 18649 12391 18683
rect 13676 18649 13710 18683
rect 17969 18649 18003 18683
rect 20370 18649 20404 18683
rect 3617 18581 3651 18615
rect 6285 18581 6319 18615
rect 8769 18581 8803 18615
rect 9965 18581 9999 18615
rect 11989 18581 12023 18615
rect 12541 18581 12575 18615
rect 15761 18581 15795 18615
rect 19257 18581 19291 18615
rect 2789 18377 2823 18411
rect 4169 18377 4203 18411
rect 4813 18377 4847 18411
rect 6009 18377 6043 18411
rect 6377 18377 6411 18411
rect 7205 18377 7239 18411
rect 8861 18377 8895 18411
rect 11253 18377 11287 18411
rect 11529 18377 11563 18411
rect 13277 18377 13311 18411
rect 14381 18377 14415 18411
rect 15025 18377 15059 18411
rect 12357 18309 12391 18343
rect 15209 18309 15243 18343
rect 17509 18309 17543 18343
rect 2973 18241 3007 18275
rect 4329 18241 4363 18275
rect 4445 18241 4479 18275
rect 4537 18241 4571 18275
rect 4721 18241 4755 18275
rect 4997 18241 5031 18275
rect 5549 18241 5583 18275
rect 6009 18241 6043 18275
rect 6193 18241 6227 18275
rect 6561 18241 6595 18275
rect 6929 18241 6963 18275
rect 7757 18241 7791 18275
rect 8309 18241 8343 18275
rect 9229 18241 9263 18275
rect 9956 18241 9990 18275
rect 11161 18241 11195 18275
rect 11345 18241 11379 18275
rect 12265 18241 12299 18275
rect 12541 18241 12575 18275
rect 12725 18241 12759 18275
rect 12909 18241 12943 18275
rect 13093 18241 13127 18275
rect 13921 18241 13955 18275
rect 14565 18241 14599 18275
rect 14924 18263 14958 18297
rect 16865 18241 16899 18275
rect 17233 18241 17267 18275
rect 17325 18241 17359 18275
rect 3249 18173 3283 18207
rect 3433 18173 3467 18207
rect 4077 18173 4111 18207
rect 5181 18173 5215 18207
rect 5641 18173 5675 18207
rect 6745 18173 6779 18207
rect 6837 18173 6871 18207
rect 7665 18173 7699 18207
rect 8401 18173 8435 18207
rect 9137 18173 9171 18207
rect 9689 18173 9723 18207
rect 12081 18173 12115 18207
rect 12817 18173 12851 18207
rect 14013 18173 14047 18207
rect 14289 18173 14323 18207
rect 14841 18173 14875 18207
rect 17141 18173 17175 18207
rect 5917 18105 5951 18139
rect 11069 18105 11103 18139
rect 15209 18105 15243 18139
rect 17509 18105 17543 18139
rect 3157 18037 3191 18071
rect 14749 18037 14783 18071
rect 16681 18037 16715 18071
rect 17049 18037 17083 18071
rect 10425 17833 10459 17867
rect 12081 17833 12115 17867
rect 14473 17833 14507 17867
rect 16129 17833 16163 17867
rect 17693 17833 17727 17867
rect 10333 17765 10367 17799
rect 4445 17697 4479 17731
rect 10977 17697 11011 17731
rect 12173 17697 12207 17731
rect 15209 17697 15243 17731
rect 15577 17697 15611 17731
rect 3433 17629 3467 17663
rect 3617 17629 3651 17663
rect 4997 17629 5031 17663
rect 9781 17629 9815 17663
rect 9965 17629 9999 17663
rect 10057 17629 10091 17663
rect 11713 17629 11747 17663
rect 11897 17629 11931 17663
rect 11989 17629 12023 17663
rect 12633 17629 12667 17663
rect 12725 17629 12759 17663
rect 13001 17629 13035 17663
rect 14657 17629 14691 17663
rect 15025 17629 15059 17663
rect 15117 17629 15151 17663
rect 15393 17629 15427 17663
rect 16037 17629 16071 17663
rect 16221 17629 16255 17663
rect 16313 17629 16347 17663
rect 16580 17629 16614 17663
rect 19717 17629 19751 17663
rect 21465 17629 21499 17663
rect 10333 17561 10367 17595
rect 11161 17561 11195 17595
rect 12817 17561 12851 17595
rect 14749 17561 14783 17595
rect 14841 17561 14875 17595
rect 3525 17493 3559 17527
rect 3801 17493 3835 17527
rect 4905 17493 4939 17527
rect 9873 17493 9907 17527
rect 10149 17493 10183 17527
rect 12449 17493 12483 17527
rect 19901 17493 19935 17527
rect 20913 17493 20947 17527
rect 3893 17289 3927 17323
rect 10701 17289 10735 17323
rect 12449 17289 12483 17323
rect 15117 17289 15151 17323
rect 21281 17289 21315 17323
rect 6377 17221 6411 17255
rect 15209 17221 15243 17255
rect 15577 17221 15611 17255
rect 20146 17221 20180 17255
rect 1409 17153 1443 17187
rect 1676 17153 1710 17187
rect 2881 17153 2915 17187
rect 3065 17153 3099 17187
rect 3617 17153 3651 17187
rect 4077 17153 4111 17187
rect 4445 17153 4479 17187
rect 4629 17153 4663 17187
rect 5641 17153 5675 17187
rect 6561 17153 6595 17187
rect 6653 17153 6687 17187
rect 7297 17153 7331 17187
rect 7481 17153 7515 17187
rect 8309 17153 8343 17187
rect 9301 17153 9335 17187
rect 12633 17153 12667 17187
rect 12817 17153 12851 17187
rect 12909 17153 12943 17187
rect 13001 17153 13035 17187
rect 13277 17153 13311 17187
rect 14473 17153 14507 17187
rect 14657 17153 14691 17187
rect 14749 17153 14783 17187
rect 14841 17153 14875 17187
rect 15393 17153 15427 17187
rect 18685 17153 18719 17187
rect 19901 17153 19935 17187
rect 3341 17085 3375 17119
rect 3801 17085 3835 17119
rect 4261 17085 4295 17119
rect 4353 17085 4387 17119
rect 8033 17085 8067 17119
rect 8125 17085 8159 17119
rect 8493 17085 8527 17119
rect 9045 17085 9079 17119
rect 11253 17085 11287 17119
rect 11621 17085 11655 17119
rect 18429 17085 18463 17119
rect 2789 17017 2823 17051
rect 7757 17017 7791 17051
rect 3249 16949 3283 16983
rect 3433 16949 3467 16983
rect 5549 16949 5583 16983
rect 6377 16949 6411 16983
rect 7481 16949 7515 16983
rect 7573 16949 7607 16983
rect 10425 16949 10459 16983
rect 12173 16949 12207 16983
rect 13093 16949 13127 16983
rect 13369 16949 13403 16983
rect 19809 16949 19843 16983
rect 3065 16745 3099 16779
rect 3433 16745 3467 16779
rect 6009 16745 6043 16779
rect 6469 16745 6503 16779
rect 12817 16745 12851 16779
rect 12909 16745 12943 16779
rect 15393 16745 15427 16779
rect 17877 16745 17911 16779
rect 19717 16745 19751 16779
rect 3249 16677 3283 16711
rect 8953 16677 8987 16711
rect 9689 16677 9723 16711
rect 11253 16677 11287 16711
rect 14933 16677 14967 16711
rect 1685 16609 1719 16643
rect 4629 16609 4663 16643
rect 7205 16609 7239 16643
rect 9873 16609 9907 16643
rect 11989 16609 12023 16643
rect 13369 16609 13403 16643
rect 15301 16609 15335 16643
rect 15761 16609 15795 16643
rect 18613 16609 18647 16643
rect 19349 16609 19383 16643
rect 19809 16609 19843 16643
rect 20361 16609 20395 16643
rect 20913 16609 20947 16643
rect 4445 16541 4479 16575
rect 6653 16541 6687 16575
rect 6929 16541 6963 16575
rect 7113 16541 7147 16575
rect 7472 16541 7506 16575
rect 9321 16541 9355 16575
rect 9505 16541 9539 16575
rect 9781 16541 9815 16575
rect 12265 16541 12299 16575
rect 12541 16541 12575 16575
rect 12633 16541 12667 16575
rect 13093 16541 13127 16575
rect 13185 16541 13219 16575
rect 13461 16541 13495 16575
rect 15577 16541 15611 16575
rect 17601 16541 17635 16575
rect 17693 16541 17727 16575
rect 18889 16541 18923 16575
rect 19073 16541 19107 16575
rect 19533 16541 19567 16575
rect 20729 16541 20763 16575
rect 21649 16541 21683 16575
rect 1952 16473 1986 16507
rect 3417 16473 3451 16507
rect 3617 16473 3651 16507
rect 4896 16473 4930 16507
rect 6745 16473 6779 16507
rect 6837 16473 6871 16507
rect 9137 16473 9171 16507
rect 10118 16473 10152 16507
rect 12449 16473 12483 16507
rect 18705 16473 18739 16507
rect 3801 16405 3835 16439
rect 8585 16405 8619 16439
rect 9781 16405 9815 16439
rect 11345 16405 11379 16439
rect 14841 16405 14875 16439
rect 17417 16405 17451 16439
rect 17969 16405 18003 16439
rect 20545 16405 20579 16439
rect 21005 16405 21039 16439
rect 3065 16201 3099 16235
rect 5733 16201 5767 16235
rect 6745 16201 6779 16235
rect 8309 16201 8343 16235
rect 11989 16201 12023 16235
rect 14657 16201 14691 16235
rect 16221 16201 16255 16235
rect 19073 16201 19107 16235
rect 19517 16201 19551 16235
rect 20177 16201 20211 16235
rect 21649 16201 21683 16235
rect 2421 16133 2455 16167
rect 4353 16133 4387 16167
rect 9597 16133 9631 16167
rect 11100 16133 11134 16167
rect 11621 16133 11655 16167
rect 12233 16133 12267 16167
rect 12449 16133 12483 16167
rect 19717 16133 19751 16167
rect 20514 16133 20548 16167
rect 2329 16065 2363 16099
rect 2513 16065 2547 16099
rect 4445 16065 4479 16099
rect 4629 16065 4663 16099
rect 4721 16065 4755 16099
rect 4813 16065 4847 16099
rect 5273 16065 5307 16099
rect 5917 16065 5951 16099
rect 6377 16065 6411 16099
rect 6561 16065 6595 16099
rect 7389 16065 7423 16099
rect 7481 16065 7515 16099
rect 7573 16065 7607 16099
rect 7757 16065 7791 16099
rect 11529 16065 11563 16099
rect 11805 16065 11839 16099
rect 12541 16065 12575 16099
rect 12725 16065 12759 16099
rect 12817 16065 12851 16099
rect 12909 16065 12943 16099
rect 14197 16065 14231 16099
rect 14381 16065 14415 16099
rect 14473 16065 14507 16099
rect 14749 16065 14783 16099
rect 15097 16065 15131 16099
rect 16957 16065 16991 16099
rect 17224 16065 17258 16099
rect 19993 16065 20027 16099
rect 5181 15997 5215 16031
rect 6193 15997 6227 16031
rect 11345 15997 11379 16031
rect 13001 15997 13035 16031
rect 14841 15997 14875 16031
rect 18429 15997 18463 16031
rect 20269 15997 20303 16031
rect 5641 15929 5675 15963
rect 6101 15929 6135 15963
rect 7113 15929 7147 15963
rect 12081 15929 12115 15963
rect 12541 15929 12575 15963
rect 14473 15929 14507 15963
rect 19349 15929 19383 15963
rect 4997 15861 5031 15895
rect 9965 15861 9999 15895
rect 12265 15861 12299 15895
rect 14381 15861 14415 15895
rect 18337 15861 18371 15895
rect 19533 15861 19567 15895
rect 2329 15657 2363 15691
rect 4537 15657 4571 15691
rect 7481 15657 7515 15691
rect 7849 15657 7883 15691
rect 13001 15657 13035 15691
rect 13277 15657 13311 15691
rect 14841 15657 14875 15691
rect 16957 15657 16991 15691
rect 18153 15657 18187 15691
rect 18797 15657 18831 15691
rect 20269 15657 20303 15691
rect 21925 15657 21959 15691
rect 2237 15521 2271 15555
rect 3801 15521 3835 15555
rect 8125 15521 8159 15555
rect 8309 15521 8343 15555
rect 19625 15521 19659 15555
rect 20085 15521 20119 15555
rect 2421 15453 2455 15487
rect 2513 15453 2547 15487
rect 2605 15453 2639 15487
rect 2697 15453 2731 15487
rect 3065 15453 3099 15487
rect 4445 15453 4479 15487
rect 4721 15453 4755 15487
rect 4997 15453 5031 15487
rect 5273 15453 5307 15487
rect 7481 15453 7515 15487
rect 7665 15453 7699 15487
rect 7757 15453 7791 15487
rect 8033 15453 8067 15487
rect 8217 15453 8251 15487
rect 13461 15453 13495 15487
rect 13645 15453 13679 15487
rect 13737 15453 13771 15487
rect 13921 15453 13955 15487
rect 14105 15453 14139 15487
rect 14657 15453 14691 15487
rect 15025 15453 15059 15487
rect 15117 15453 15151 15487
rect 15209 15453 15243 15487
rect 15301 15453 15335 15487
rect 15669 15453 15703 15487
rect 17509 15453 17543 15487
rect 18245 15453 18279 15487
rect 18429 15453 18463 15487
rect 19073 15453 19107 15487
rect 19441 15453 19475 15487
rect 19993 15453 20027 15487
rect 20545 15453 20579 15487
rect 2881 15385 2915 15419
rect 5181 15385 5215 15419
rect 13185 15385 13219 15419
rect 19257 15385 19291 15419
rect 20269 15385 20303 15419
rect 20812 15385 20846 15419
rect 2605 15317 2639 15351
rect 3617 15317 3651 15351
rect 4905 15317 4939 15351
rect 12817 15317 12851 15351
rect 12985 15317 13019 15351
rect 13829 15317 13863 15351
rect 18521 15317 18555 15351
rect 18613 15317 18647 15351
rect 18889 15317 18923 15351
rect 19809 15317 19843 15351
rect 2789 15113 2823 15147
rect 4721 15113 4755 15147
rect 13829 15113 13863 15147
rect 14749 15113 14783 15147
rect 15485 15113 15519 15147
rect 16681 15113 16715 15147
rect 19809 15113 19843 15147
rect 20913 15113 20947 15147
rect 1676 15045 1710 15079
rect 3157 15045 3191 15079
rect 3373 15045 3407 15079
rect 4813 15045 4847 15079
rect 6469 15045 6503 15079
rect 18245 15045 18279 15079
rect 19961 15045 19995 15079
rect 20177 15045 20211 15079
rect 1409 14977 1443 15011
rect 3801 14977 3835 15011
rect 4169 14977 4203 15011
rect 4445 14977 4479 15011
rect 4537 14977 4571 15011
rect 4997 14977 5031 15011
rect 5089 14977 5123 15011
rect 12173 14977 12207 15011
rect 12449 14977 12483 15011
rect 12705 14977 12739 15011
rect 14289 14977 14323 15011
rect 14565 14977 14599 15011
rect 15577 14977 15611 15011
rect 17805 14977 17839 15011
rect 18061 14977 18095 15011
rect 18429 14977 18463 15011
rect 18521 14977 18555 15011
rect 18797 14977 18831 15011
rect 19073 14977 19107 15011
rect 19257 14977 19291 15011
rect 19533 14977 19567 15011
rect 20269 14977 20303 15011
rect 20453 14977 20487 15011
rect 20637 14977 20671 15011
rect 20729 14977 20763 15011
rect 3617 14909 3651 14943
rect 4077 14909 4111 14943
rect 4261 14909 4295 14943
rect 3525 14841 3559 14875
rect 4813 14841 4847 14875
rect 12357 14841 12391 14875
rect 18705 14841 18739 14875
rect 18981 14841 19015 14875
rect 3341 14773 3375 14807
rect 3985 14773 4019 14807
rect 6745 14773 6779 14807
rect 14381 14773 14415 14807
rect 18429 14773 18463 14807
rect 19717 14773 19751 14807
rect 19993 14773 20027 14807
rect 3433 14569 3467 14603
rect 3893 14569 3927 14603
rect 5365 14569 5399 14603
rect 7849 14569 7883 14603
rect 9689 14569 9723 14603
rect 13001 14569 13035 14603
rect 14565 14569 14599 14603
rect 14749 14569 14783 14603
rect 15209 14569 15243 14603
rect 18429 14569 18463 14603
rect 6009 14501 6043 14535
rect 8677 14501 8711 14535
rect 9137 14501 9171 14535
rect 13185 14501 13219 14535
rect 2053 14433 2087 14467
rect 4445 14433 4479 14467
rect 8953 14433 8987 14467
rect 15393 14433 15427 14467
rect 15669 14433 15703 14467
rect 16589 14433 16623 14467
rect 17049 14433 17083 14467
rect 19257 14433 19291 14467
rect 2320 14365 2354 14399
rect 5181 14365 5215 14399
rect 5549 14365 5583 14399
rect 5641 14365 5675 14399
rect 5825 14365 5859 14399
rect 5917 14365 5951 14399
rect 6193 14365 6227 14399
rect 6285 14365 6319 14399
rect 6745 14365 6779 14399
rect 7021 14365 7055 14399
rect 7113 14365 7147 14399
rect 7481 14365 7515 14399
rect 7665 14365 7699 14399
rect 8033 14365 8067 14399
rect 8309 14365 8343 14399
rect 8493 14365 8527 14399
rect 8585 14365 8619 14399
rect 9505 14365 9539 14399
rect 9873 14365 9907 14399
rect 10057 14365 10091 14399
rect 10701 14365 10735 14399
rect 11161 14365 11195 14399
rect 12817 14365 12851 14399
rect 13093 14365 13127 14399
rect 13369 14365 13403 14399
rect 13461 14365 13495 14399
rect 15117 14365 15151 14399
rect 15485 14365 15519 14399
rect 15577 14365 15611 14399
rect 16773 14365 16807 14399
rect 19533 14365 19567 14399
rect 4629 14297 4663 14331
rect 6009 14297 6043 14331
rect 6561 14297 6595 14331
rect 6929 14297 6963 14331
rect 7205 14297 7239 14331
rect 9413 14297 9447 14331
rect 13185 14297 13219 14331
rect 14749 14297 14783 14331
rect 17316 14297 17350 14331
rect 7481 14229 7515 14263
rect 9965 14229 9999 14263
rect 10885 14229 10919 14263
rect 11345 14229 11379 14263
rect 12633 14229 12667 14263
rect 16957 14229 16991 14263
rect 20269 14229 20303 14263
rect 5279 14025 5313 14059
rect 5365 14025 5399 14059
rect 8493 14025 8527 14059
rect 9965 14025 9999 14059
rect 11529 14025 11563 14059
rect 13461 14025 13495 14059
rect 14381 14025 14415 14059
rect 15393 14025 15427 14059
rect 16037 14025 16071 14059
rect 17509 14025 17543 14059
rect 8585 13957 8619 13991
rect 9873 13957 9907 13991
rect 11078 13957 11112 13991
rect 12326 13957 12360 13991
rect 16189 13957 16223 13991
rect 16405 13957 16439 13991
rect 3157 13889 3191 13923
rect 3341 13889 3375 13923
rect 3433 13889 3467 13923
rect 3689 13889 3723 13923
rect 5181 13889 5215 13923
rect 5457 13889 5491 13923
rect 5733 13889 5767 13923
rect 6561 13889 6595 13923
rect 6653 13889 6687 13923
rect 6745 13889 6779 13923
rect 7113 13889 7147 13923
rect 7380 13889 7414 13923
rect 8861 13889 8895 13923
rect 9321 13889 9355 13923
rect 11713 13889 11747 13923
rect 11897 13889 11931 13923
rect 14841 13889 14875 13923
rect 15485 13889 15519 13923
rect 17325 13889 17359 13923
rect 17785 13889 17819 13923
rect 18521 13889 18555 13923
rect 19993 13889 20027 13923
rect 20260 13889 20294 13923
rect 3249 13821 3283 13855
rect 5825 13821 5859 13855
rect 6837 13821 6871 13855
rect 11345 13821 11379 13855
rect 12081 13821 12115 13855
rect 14933 13821 14967 13855
rect 15945 13821 15979 13855
rect 17141 13821 17175 13855
rect 17877 13821 17911 13855
rect 4813 13753 4847 13787
rect 6101 13753 6135 13787
rect 8953 13753 8987 13787
rect 9045 13753 9079 13787
rect 9413 13753 9447 13787
rect 9597 13753 9631 13787
rect 15209 13753 15243 13787
rect 17601 13753 17635 13787
rect 7021 13685 7055 13719
rect 9137 13685 9171 13719
rect 14565 13685 14599 13719
rect 15669 13685 15703 13719
rect 16221 13685 16255 13719
rect 21373 13685 21407 13719
rect 8493 13481 8527 13515
rect 9413 13481 9447 13515
rect 10517 13481 10551 13515
rect 15393 13481 15427 13515
rect 15669 13481 15703 13515
rect 9321 13413 9355 13447
rect 9689 13413 9723 13447
rect 13553 13413 13587 13447
rect 15209 13413 15243 13447
rect 5365 13345 5399 13379
rect 8953 13345 8987 13379
rect 10241 13345 10275 13379
rect 11069 13345 11103 13379
rect 12173 13345 12207 13379
rect 14565 13345 14599 13379
rect 20545 13345 20579 13379
rect 5632 13277 5666 13311
rect 7021 13277 7055 13311
rect 7849 13277 7883 13311
rect 8217 13277 8251 13311
rect 8309 13277 8343 13311
rect 10057 13277 10091 13311
rect 10977 13277 11011 13311
rect 15301 13277 15335 13311
rect 15485 13277 15519 13311
rect 17049 13277 17083 13311
rect 18705 13277 18739 13311
rect 18797 13277 18831 13311
rect 18981 13277 19015 13311
rect 19441 13277 19475 13311
rect 19533 13277 19567 13311
rect 20453 13277 20487 13311
rect 20729 13277 20763 13311
rect 20913 13277 20947 13311
rect 21005 13277 21039 13311
rect 21557 13277 21591 13311
rect 8033 13209 8067 13243
rect 10885 13209 10919 13243
rect 12418 13209 12452 13243
rect 16782 13209 16816 13243
rect 6745 13141 6779 13175
rect 7205 13141 7239 13175
rect 10149 13141 10183 13175
rect 14749 13141 14783 13175
rect 14841 13141 14875 13175
rect 19257 13141 19291 13175
rect 19717 13141 19751 13175
rect 19809 13141 19843 13175
rect 7297 12937 7331 12971
rect 13001 12937 13035 12971
rect 16497 12937 16531 12971
rect 19717 12937 19751 12971
rect 21465 12937 21499 12971
rect 6837 12869 6871 12903
rect 11713 12869 11747 12903
rect 18245 12869 18279 12903
rect 3709 12801 3743 12835
rect 7021 12801 7055 12835
rect 7113 12801 7147 12835
rect 7205 12801 7239 12835
rect 7389 12801 7423 12835
rect 15301 12801 15335 12835
rect 16037 12801 16071 12835
rect 16221 12801 16255 12835
rect 16313 12801 16347 12835
rect 17969 12801 18003 12835
rect 18153 12801 18187 12835
rect 20085 12801 20119 12835
rect 20341 12801 20375 12835
rect 3525 12733 3559 12767
rect 15393 12733 15427 12767
rect 15577 12733 15611 12767
rect 15853 12733 15887 12767
rect 6837 12665 6871 12699
rect 14933 12665 14967 12699
rect 3893 12597 3927 12631
rect 17785 12597 17819 12631
rect 3801 12393 3835 12427
rect 10517 12393 10551 12427
rect 11989 12393 12023 12427
rect 21465 12393 21499 12427
rect 3433 12325 3467 12359
rect 19257 12325 19291 12359
rect 4353 12257 4387 12291
rect 17601 12257 17635 12291
rect 2053 12189 2087 12223
rect 4721 12189 4755 12223
rect 5273 12189 5307 12223
rect 5549 12189 5583 12223
rect 5733 12189 5767 12223
rect 5917 12189 5951 12223
rect 6193 12189 6227 12223
rect 9137 12189 9171 12223
rect 10885 12189 10919 12223
rect 11069 12189 11103 12223
rect 11253 12189 11287 12223
rect 11805 12189 11839 12223
rect 14473 12189 14507 12223
rect 17325 12189 17359 12223
rect 19809 12189 19843 12223
rect 20177 12189 20211 12223
rect 20361 12189 20395 12223
rect 20453 12189 20487 12223
rect 20729 12189 20763 12223
rect 2298 12121 2332 12155
rect 9404 12121 9438 12155
rect 17846 12121 17880 12155
rect 4537 12053 4571 12087
rect 5089 12053 5123 12087
rect 6009 12053 6043 12087
rect 14289 12053 14323 12087
rect 17509 12053 17543 12087
rect 18981 12053 19015 12087
rect 19993 12053 20027 12087
rect 5549 11849 5583 11883
rect 8677 11849 8711 11883
rect 10333 11849 10367 11883
rect 15577 11849 15611 11883
rect 20177 11849 20211 11883
rect 21097 11849 21131 11883
rect 4344 11781 4378 11815
rect 6377 11781 6411 11815
rect 6593 11781 6627 11815
rect 9413 11781 9447 11815
rect 15945 11781 15979 11815
rect 18328 11781 18362 11815
rect 21005 11781 21039 11815
rect 1501 11713 1535 11747
rect 1768 11713 1802 11747
rect 4077 11713 4111 11747
rect 6929 11713 6963 11747
rect 7113 11713 7147 11747
rect 7389 11713 7423 11747
rect 7941 11713 7975 11747
rect 9965 11713 9999 11747
rect 10057 11713 10091 11747
rect 10241 11713 10275 11747
rect 10517 11713 10551 11747
rect 10793 11713 10827 11747
rect 11345 11713 11379 11747
rect 12541 11713 12575 11747
rect 12909 11713 12943 11747
rect 13093 11713 13127 11747
rect 13369 11713 13403 11747
rect 13921 11713 13955 11747
rect 15209 11713 15243 11747
rect 15669 11713 15703 11747
rect 15853 11713 15887 11747
rect 16313 11713 16347 11747
rect 18061 11713 18095 11747
rect 20361 11713 20395 11747
rect 20545 11713 20579 11747
rect 20821 11713 20855 11747
rect 21281 11713 21315 11747
rect 21649 11713 21683 11747
rect 3709 11645 3743 11679
rect 6193 11645 6227 11679
rect 7573 11645 7607 11679
rect 7665 11645 7699 11679
rect 10977 11645 11011 11679
rect 12265 11645 12299 11679
rect 13553 11645 13587 11679
rect 13645 11645 13679 11679
rect 14933 11645 14967 11679
rect 16129 11645 16163 11679
rect 16681 11645 16715 11679
rect 17233 11645 17267 11679
rect 19625 11645 19659 11679
rect 2881 11577 2915 11611
rect 9689 11577 9723 11611
rect 14657 11577 14691 11611
rect 21465 11577 21499 11611
rect 3157 11509 3191 11543
rect 5457 11509 5491 11543
rect 6561 11509 6595 11543
rect 6745 11509 6779 11543
rect 10609 11509 10643 11543
rect 11161 11509 11195 11543
rect 11621 11509 11655 11543
rect 12357 11509 12391 11543
rect 16497 11509 16531 11543
rect 19441 11509 19475 11543
rect 1685 11305 1719 11339
rect 2145 11305 2179 11339
rect 3433 11305 3467 11339
rect 4353 11305 4387 11339
rect 9781 11305 9815 11339
rect 11805 11305 11839 11339
rect 13921 11305 13955 11339
rect 14473 11305 14507 11339
rect 14749 11305 14783 11339
rect 15209 11305 15243 11339
rect 16037 11305 16071 11339
rect 19257 11305 19291 11339
rect 19717 11305 19751 11339
rect 20361 11305 20395 11339
rect 20637 11305 20671 11339
rect 20821 11305 20855 11339
rect 3617 11237 3651 11271
rect 7113 11237 7147 11271
rect 9229 11237 9263 11271
rect 13277 11237 13311 11271
rect 13369 11237 13403 11271
rect 14289 11237 14323 11271
rect 19073 11237 19107 11271
rect 2237 11169 2271 11203
rect 3065 11169 3099 11203
rect 4629 11169 4663 11203
rect 17417 11169 17451 11203
rect 19809 11169 19843 11203
rect 1869 11101 1903 11135
rect 1961 11101 1995 11135
rect 2421 11101 2455 11135
rect 2605 11101 2639 11135
rect 2881 11101 2915 11135
rect 3341 11101 3375 11135
rect 3433 11101 3467 11135
rect 3985 11101 4019 11135
rect 4077 11101 4111 11135
rect 4896 11101 4930 11135
rect 6377 11101 6411 11135
rect 8493 11101 8527 11135
rect 10333 11101 10367 11135
rect 10425 11101 10459 11135
rect 11897 11101 11931 11135
rect 14933 11101 14967 11135
rect 15025 11101 15059 11135
rect 15301 11101 15335 11135
rect 18889 11101 18923 11135
rect 19441 11101 19475 11135
rect 19533 11101 19567 11135
rect 20085 11101 20119 11135
rect 20177 11101 20211 11135
rect 2697 11033 2731 11067
rect 3157 11033 3191 11067
rect 3801 11033 3835 11067
rect 4169 11033 4203 11067
rect 8226 11033 8260 11067
rect 9045 11033 9079 11067
rect 9689 11033 9723 11067
rect 10692 11033 10726 11067
rect 12164 11033 12198 11067
rect 14457 11033 14491 11067
rect 14657 11033 14691 11067
rect 15209 11033 15243 11067
rect 17150 11033 17184 11067
rect 19717 11033 19751 11067
rect 20453 11033 20487 11067
rect 20653 11033 20687 11067
rect 6009 10965 6043 10999
rect 7021 10965 7055 10999
rect 10149 10965 10183 10999
rect 13553 10965 13587 10999
rect 13645 10965 13679 10999
rect 13737 10965 13771 10999
rect 15945 10965 15979 10999
rect 19993 10965 20027 10999
rect 3341 10761 3375 10795
rect 6193 10761 6227 10795
rect 7021 10761 7055 10795
rect 7757 10761 7791 10795
rect 8033 10761 8067 10795
rect 11529 10761 11563 10795
rect 12817 10761 12851 10795
rect 15301 10761 15335 10795
rect 16865 10761 16899 10795
rect 16957 10761 16991 10795
rect 5080 10693 5114 10727
rect 10232 10693 10266 10727
rect 15669 10693 15703 10727
rect 18070 10693 18104 10727
rect 19778 10693 19812 10727
rect 15439 10659 15473 10693
rect 2329 10625 2363 10659
rect 3893 10625 3927 10659
rect 4813 10625 4847 10659
rect 6561 10625 6595 10659
rect 6837 10625 6871 10659
rect 7113 10625 7147 10659
rect 7297 10625 7331 10659
rect 7481 10625 7515 10659
rect 7573 10625 7607 10659
rect 7849 10625 7883 10659
rect 11713 10625 11747 10659
rect 11805 10625 11839 10659
rect 12633 10625 12667 10659
rect 13829 10625 13863 10659
rect 14096 10625 14130 10659
rect 15945 10625 15979 10659
rect 16037 10625 16071 10659
rect 16313 10625 16347 10659
rect 16681 10625 16715 10659
rect 18337 10625 18371 10659
rect 19533 10625 19567 10659
rect 2513 10557 2547 10591
rect 2605 10557 2639 10591
rect 3157 10557 3191 10591
rect 6653 10557 6687 10591
rect 9965 10557 9999 10591
rect 13461 10557 13495 10591
rect 21005 10557 21039 10591
rect 11345 10489 11379 10523
rect 2145 10421 2179 10455
rect 6653 10421 6687 10455
rect 12081 10421 12115 10455
rect 15209 10421 15243 10455
rect 15485 10421 15519 10455
rect 15761 10421 15795 10455
rect 16497 10421 16531 10455
rect 20913 10421 20947 10455
rect 21649 10421 21683 10455
rect 3525 10217 3559 10251
rect 4997 10217 5031 10251
rect 6561 10217 6595 10251
rect 6745 10217 6779 10251
rect 12541 10217 12575 10251
rect 13369 10217 13403 10251
rect 14841 10217 14875 10251
rect 20637 10217 20671 10251
rect 20729 10217 20763 10251
rect 20913 10217 20947 10251
rect 13553 10149 13587 10183
rect 16865 10149 16899 10183
rect 2145 10081 2179 10115
rect 6009 10081 6043 10115
rect 12173 10081 12207 10115
rect 13277 10081 13311 10115
rect 14657 10081 14691 10115
rect 17693 10081 17727 10115
rect 21649 10081 21683 10115
rect 1869 10013 1903 10047
rect 5181 10013 5215 10047
rect 5365 10013 5399 10047
rect 5457 10013 5491 10047
rect 9229 10013 9263 10047
rect 9413 10013 9447 10047
rect 12357 10013 12391 10047
rect 13369 10013 13403 10047
rect 15025 10013 15059 10047
rect 15209 10013 15243 10047
rect 15485 10013 15519 10047
rect 19073 10013 19107 10047
rect 19257 10013 19291 10047
rect 20913 10013 20947 10047
rect 21005 10013 21039 10047
rect 21465 10013 21499 10047
rect 2390 9945 2424 9979
rect 6377 9945 6411 9979
rect 6577 9945 6611 9979
rect 13093 9945 13127 9979
rect 15730 9945 15764 9979
rect 19502 9945 19536 9979
rect 21189 9945 21223 9979
rect 2053 9877 2087 9911
rect 9321 9877 9355 9911
rect 14105 9877 14139 9911
rect 15393 9877 15427 9911
rect 17141 9877 17175 9911
rect 18429 9877 18463 9911
rect 21281 9877 21315 9911
rect 2973 9673 3007 9707
rect 9873 9673 9907 9707
rect 16957 9673 16991 9707
rect 19165 9673 19199 9707
rect 20805 9673 20839 9707
rect 8033 9605 8067 9639
rect 9514 9605 9548 9639
rect 13737 9605 13771 9639
rect 21005 9605 21039 9639
rect 1593 9537 1627 9571
rect 1860 9537 1894 9571
rect 3985 9537 4019 9571
rect 4169 9537 4203 9571
rect 5457 9537 5491 9571
rect 5825 9537 5859 9571
rect 5917 9537 5951 9571
rect 6101 9537 6135 9571
rect 7297 9537 7331 9571
rect 8217 9537 8251 9571
rect 8309 9537 8343 9571
rect 10149 9537 10183 9571
rect 11621 9537 11655 9571
rect 11805 9537 11839 9571
rect 13553 9537 13587 9571
rect 17141 9537 17175 9571
rect 18429 9537 18463 9571
rect 18613 9537 18647 9571
rect 18797 9537 18831 9571
rect 18889 9537 18923 9571
rect 20289 9537 20323 9571
rect 21281 9537 21315 9571
rect 5733 9469 5767 9503
rect 9781 9469 9815 9503
rect 10058 9469 10092 9503
rect 10241 9469 10275 9503
rect 10333 9469 10367 9503
rect 13369 9469 13403 9503
rect 17325 9469 17359 9503
rect 20545 9469 20579 9503
rect 19073 9401 19107 9435
rect 20637 9401 20671 9435
rect 3985 9333 4019 9367
rect 5273 9333 5307 9367
rect 5641 9333 5675 9367
rect 6101 9333 6135 9367
rect 7205 9333 7239 9367
rect 8033 9333 8067 9367
rect 8401 9333 8435 9367
rect 11805 9333 11839 9367
rect 20821 9333 20855 9367
rect 21097 9333 21131 9367
rect 2237 9129 2271 9163
rect 4353 9129 4387 9163
rect 5917 9129 5951 9163
rect 8585 9129 8619 9163
rect 8953 9129 8987 9163
rect 11805 9129 11839 9163
rect 11897 9129 11931 9163
rect 14105 9129 14139 9163
rect 20453 9129 20487 9163
rect 21925 9129 21959 9163
rect 1593 9061 1627 9095
rect 9965 9061 9999 9095
rect 10241 9061 10275 9095
rect 3985 8993 4019 9027
rect 5181 8993 5215 9027
rect 5825 8993 5859 9027
rect 11345 8993 11379 9027
rect 11437 8993 11471 9027
rect 20545 8993 20579 9027
rect 1409 8925 1443 8959
rect 1869 8925 1903 8959
rect 1961 8925 1995 8959
rect 2145 8925 2179 8959
rect 2421 8925 2455 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 4997 8925 5031 8959
rect 6561 8925 6595 8959
rect 8125 8925 8159 8959
rect 8401 8925 8435 8959
rect 8677 8925 8711 8959
rect 9229 8925 9263 8959
rect 9321 8925 9355 8959
rect 9413 8925 9447 8959
rect 9597 8925 9631 8959
rect 10885 8925 10919 8959
rect 11069 8925 11103 8959
rect 11161 8925 11195 8959
rect 11529 8925 11563 8959
rect 11621 8925 11655 8959
rect 12081 8925 12115 8959
rect 12357 8925 12391 8959
rect 12541 8925 12575 8959
rect 12817 8925 12851 8959
rect 15485 8925 15519 8959
rect 17233 8925 17267 8959
rect 17417 8925 17451 8959
rect 19901 8925 19935 8959
rect 19993 8925 20027 8959
rect 20177 8925 20211 8959
rect 20269 8925 20303 8959
rect 20812 8925 20846 8959
rect 7880 8857 7914 8891
rect 9689 8857 9723 8891
rect 10425 8857 10459 8891
rect 10609 8857 10643 8891
rect 15218 8857 15252 8891
rect 4261 8789 4295 8823
rect 6745 8789 6779 8823
rect 8217 8789 8251 8823
rect 10149 8789 10183 8823
rect 10701 8789 10735 8823
rect 12725 8789 12759 8823
rect 17049 8789 17083 8823
rect 6101 8585 6135 8619
rect 6377 8585 6411 8619
rect 9505 8585 9539 8619
rect 10057 8585 10091 8619
rect 10510 8585 10544 8619
rect 11345 8585 11379 8619
rect 12909 8585 12943 8619
rect 16037 8585 16071 8619
rect 16497 8585 16531 8619
rect 18153 8585 18187 8619
rect 20913 8585 20947 8619
rect 3424 8517 3458 8551
rect 4988 8517 5022 8551
rect 8125 8517 8159 8551
rect 9137 8517 9171 8551
rect 10241 8517 10275 8551
rect 16926 8517 16960 8551
rect 7573 8449 7607 8483
rect 8033 8449 8067 8483
rect 8309 8449 8343 8483
rect 8953 8449 8987 8483
rect 9045 8449 9079 8483
rect 9229 8449 9263 8483
rect 9413 8449 9447 8483
rect 9689 8449 9723 8483
rect 9965 8449 9999 8483
rect 10333 8449 10367 8483
rect 10425 8449 10459 8483
rect 10609 8449 10643 8483
rect 11785 8449 11819 8483
rect 13645 8449 13679 8483
rect 13737 8449 13771 8483
rect 14269 8449 14303 8483
rect 15853 8449 15887 8483
rect 16313 8449 16347 8483
rect 16681 8449 16715 8483
rect 21465 8449 21499 8483
rect 3157 8381 3191 8415
rect 4721 8381 4755 8415
rect 6929 8381 6963 8415
rect 7481 8381 7515 8415
rect 9873 8381 9907 8415
rect 10793 8381 10827 8415
rect 11529 8381 11563 8415
rect 14013 8381 14047 8415
rect 18705 8381 18739 8415
rect 7941 8313 7975 8347
rect 8493 8313 8527 8347
rect 8769 8313 8803 8347
rect 13461 8313 13495 8347
rect 4537 8245 4571 8279
rect 10241 8245 10275 8279
rect 13829 8245 13863 8279
rect 15393 8245 15427 8279
rect 18061 8245 18095 8279
rect 7665 8041 7699 8075
rect 8033 8041 8067 8075
rect 8585 8041 8619 8075
rect 10149 8041 10183 8075
rect 12081 8041 12115 8075
rect 13921 8041 13955 8075
rect 14749 8041 14783 8075
rect 17693 8041 17727 8075
rect 11897 7973 11931 8007
rect 7205 7905 7239 7939
rect 8217 7905 8251 7939
rect 16313 7905 16347 7939
rect 18061 7905 18095 7939
rect 21097 7905 21131 7939
rect 21557 7905 21591 7939
rect 3801 7837 3835 7871
rect 5273 7837 5307 7871
rect 7113 7837 7147 7871
rect 7389 7837 7423 7871
rect 7481 7837 7515 7871
rect 7757 7837 7791 7871
rect 8401 7837 8435 7871
rect 9873 7837 9907 7871
rect 10149 7837 10183 7871
rect 10517 7837 10551 7871
rect 12357 7837 12391 7871
rect 12449 7837 12483 7871
rect 12541 7837 12575 7871
rect 12633 7837 12667 7871
rect 12817 7837 12851 7871
rect 13737 7837 13771 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 14473 7837 14507 7871
rect 14565 7837 14599 7871
rect 15117 7837 15151 7871
rect 15301 7837 15335 7871
rect 15485 7837 15519 7871
rect 16037 7837 16071 7871
rect 19441 7837 19475 7871
rect 20177 7837 20211 7871
rect 20545 7837 20579 7871
rect 21373 7837 21407 7871
rect 21833 7837 21867 7871
rect 4068 7769 4102 7803
rect 8043 7769 8077 7803
rect 10762 7769 10796 7803
rect 16558 7769 16592 7803
rect 21189 7769 21223 7803
rect 5181 7701 5215 7735
rect 6561 7701 6595 7735
rect 7849 7701 7883 7735
rect 9965 7701 9999 7735
rect 16221 7701 16255 7735
rect 18705 7701 18739 7735
rect 19257 7701 19291 7735
rect 20361 7701 20395 7735
rect 21649 7701 21683 7735
rect 5575 7497 5609 7531
rect 6469 7497 6503 7531
rect 11529 7497 11563 7531
rect 13921 7497 13955 7531
rect 19533 7497 19567 7531
rect 20269 7497 20303 7531
rect 4353 7429 4387 7463
rect 5365 7429 5399 7463
rect 8033 7429 8067 7463
rect 14565 7429 14599 7463
rect 6653 7361 6687 7395
rect 6745 7361 6779 7395
rect 6929 7361 6963 7395
rect 7031 7351 7065 7385
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 7481 7361 7515 7395
rect 7665 7361 7699 7395
rect 8125 7361 8159 7395
rect 11897 7361 11931 7395
rect 13829 7361 13863 7395
rect 14013 7361 14047 7395
rect 14473 7361 14507 7395
rect 17785 7361 17819 7395
rect 17969 7361 18003 7395
rect 18245 7361 18279 7395
rect 18797 7361 18831 7395
rect 19809 7361 19843 7395
rect 20085 7361 20119 7395
rect 21393 7361 21427 7395
rect 21649 7361 21683 7395
rect 11989 7293 12023 7327
rect 14749 7293 14783 7327
rect 17509 7293 17543 7327
rect 18429 7293 18463 7327
rect 18521 7293 18555 7327
rect 19901 7293 19935 7327
rect 7113 7225 7147 7259
rect 19625 7225 19659 7259
rect 3065 7157 3099 7191
rect 5549 7157 5583 7191
rect 5733 7157 5767 7191
rect 14105 7157 14139 7191
rect 16865 7157 16899 7191
rect 20085 7157 20119 7191
rect 13461 6953 13495 6987
rect 16681 6953 16715 6987
rect 17969 6953 18003 6987
rect 18245 6953 18279 6987
rect 19257 6953 19291 6987
rect 19441 6953 19475 6987
rect 19901 6953 19935 6987
rect 9597 6885 9631 6919
rect 13645 6885 13679 6919
rect 17693 6885 17727 6919
rect 4813 6817 4847 6851
rect 10057 6817 10091 6851
rect 10720 6817 10754 6851
rect 11989 6817 12023 6851
rect 14657 6817 14691 6851
rect 17141 6817 17175 6851
rect 17877 6817 17911 6851
rect 20545 6817 20579 6851
rect 5089 6749 5123 6783
rect 5273 6749 5307 6783
rect 8033 6749 8067 6783
rect 8309 6749 8343 6783
rect 9045 6749 9079 6783
rect 9229 6749 9263 6783
rect 9505 6749 9539 6783
rect 9965 6749 9999 6783
rect 10241 6749 10275 6783
rect 10425 6749 10459 6783
rect 10517 6749 10551 6783
rect 11713 6749 11747 6783
rect 11897 6749 11931 6783
rect 14473 6749 14507 6783
rect 15117 6749 15151 6783
rect 15301 6749 15335 6783
rect 16313 6749 16347 6783
rect 16865 6749 16899 6783
rect 16957 6749 16991 6783
rect 17325 6749 17359 6783
rect 18061 6749 18095 6783
rect 18429 6749 18463 6783
rect 18521 6749 18555 6783
rect 18705 6749 18739 6783
rect 18981 6749 19015 6783
rect 20812 6749 20846 6783
rect 8217 6681 8251 6715
rect 9873 6681 9907 6715
rect 10793 6681 10827 6715
rect 13921 6681 13955 6715
rect 17785 6681 17819 6715
rect 19625 6681 19659 6715
rect 20085 6681 20119 6715
rect 4169 6613 4203 6647
rect 4905 6613 4939 6647
rect 8131 6613 8165 6647
rect 10609 6613 10643 6647
rect 14105 6613 14139 6647
rect 14565 6613 14599 6647
rect 15485 6613 15519 6647
rect 16497 6613 16531 6647
rect 17417 6613 17451 6647
rect 17509 6613 17543 6647
rect 18797 6613 18831 6647
rect 19425 6613 19459 6647
rect 19717 6613 19751 6647
rect 19885 6613 19919 6647
rect 21925 6613 21959 6647
rect 9229 6409 9263 6443
rect 9873 6409 9907 6443
rect 11713 6409 11747 6443
rect 13185 6409 13219 6443
rect 13921 6409 13955 6443
rect 15393 6409 15427 6443
rect 18061 6409 18095 6443
rect 19533 6409 19567 6443
rect 5304 6341 5338 6375
rect 5733 6341 5767 6375
rect 8217 6341 8251 6375
rect 10232 6341 10266 6375
rect 12357 6341 12391 6375
rect 12633 6341 12667 6375
rect 13645 6341 13679 6375
rect 15056 6341 15090 6375
rect 3985 6273 4019 6307
rect 4077 6273 4111 6307
rect 5641 6273 5675 6307
rect 5825 6273 5859 6307
rect 6561 6273 6595 6307
rect 6745 6273 6779 6307
rect 6837 6273 6871 6307
rect 7113 6273 7147 6307
rect 7757 6273 7791 6307
rect 8401 6273 8435 6307
rect 8585 6273 8619 6307
rect 8677 6273 8711 6307
rect 8861 6273 8895 6307
rect 9045 6273 9079 6307
rect 9505 6273 9539 6307
rect 11897 6273 11931 6307
rect 11989 6273 12023 6307
rect 12173 6273 12207 6307
rect 15577 6273 15611 6307
rect 16681 6273 16715 6307
rect 16937 6273 16971 6307
rect 18153 6273 18187 6307
rect 18420 6273 18454 6307
rect 19625 6273 19659 6307
rect 19892 6273 19926 6307
rect 3801 6205 3835 6239
rect 5549 6205 5583 6239
rect 6929 6205 6963 6239
rect 7849 6205 7883 6239
rect 9597 6205 9631 6239
rect 9965 6205 9999 6239
rect 15301 6205 15335 6239
rect 15853 6205 15887 6239
rect 3893 6137 3927 6171
rect 8125 6137 8159 6171
rect 13001 6137 13035 6171
rect 13277 6137 13311 6171
rect 4169 6069 4203 6103
rect 7297 6069 7331 6103
rect 11345 6069 11379 6103
rect 13093 6069 13127 6103
rect 16497 6069 16531 6103
rect 21005 6069 21039 6103
rect 6469 5865 6503 5899
rect 6929 5865 6963 5899
rect 8677 5865 8711 5899
rect 9781 5865 9815 5899
rect 15485 5865 15519 5899
rect 16037 5865 16071 5899
rect 20269 5865 20303 5899
rect 5457 5797 5491 5831
rect 6285 5797 6319 5831
rect 9413 5729 9447 5763
rect 10609 5729 10643 5763
rect 11253 5729 11287 5763
rect 16497 5729 16531 5763
rect 19625 5729 19659 5763
rect 21189 5729 21223 5763
rect 4077 5661 4111 5695
rect 6101 5661 6135 5695
rect 8309 5661 8343 5695
rect 8585 5661 8619 5695
rect 8769 5661 8803 5695
rect 9597 5661 9631 5695
rect 9873 5661 9907 5695
rect 10425 5661 10459 5695
rect 10701 5661 10735 5695
rect 11161 5661 11195 5695
rect 11805 5661 11839 5695
rect 12909 5661 12943 5695
rect 14105 5661 14139 5695
rect 15853 5661 15887 5695
rect 16129 5661 16163 5695
rect 16313 5661 16347 5695
rect 18613 5661 18647 5695
rect 20453 5661 20487 5695
rect 4344 5593 4378 5627
rect 6453 5593 6487 5627
rect 6653 5593 6687 5627
rect 8064 5593 8098 5627
rect 12173 5593 12207 5627
rect 14350 5593 14384 5627
rect 5549 5525 5583 5559
rect 12725 5525 12759 5559
rect 18061 5525 18095 5559
rect 20177 5525 20211 5559
rect 20637 5525 20671 5559
rect 4537 5321 4571 5355
rect 9873 5321 9907 5355
rect 15301 5321 15335 5355
rect 19717 5321 19751 5355
rect 20453 5321 20487 5355
rect 20913 5321 20947 5355
rect 5181 5253 5215 5287
rect 7757 5253 7791 5287
rect 14749 5253 14783 5287
rect 18245 5253 18279 5287
rect 4721 5185 4755 5219
rect 4905 5185 4939 5219
rect 5089 5185 5123 5219
rect 5273 5185 5307 5219
rect 7021 5185 7055 5219
rect 7205 5185 7239 5219
rect 7297 5185 7331 5219
rect 7389 5185 7423 5219
rect 7849 5185 7883 5219
rect 8401 5185 8435 5219
rect 9781 5185 9815 5219
rect 9965 5185 9999 5219
rect 16037 5185 16071 5219
rect 17785 5185 17819 5219
rect 17969 5185 18003 5219
rect 20085 5185 20119 5219
rect 20269 5185 20303 5219
rect 20637 5185 20671 5219
rect 20729 5185 20763 5219
rect 4997 5117 5031 5151
rect 8309 5117 8343 5151
rect 16313 5117 16347 5151
rect 7573 4981 7607 5015
rect 13277 4981 13311 5015
rect 17601 4981 17635 5015
rect 13829 4777 13863 4811
rect 16129 4777 16163 4811
rect 16221 4709 16255 4743
rect 7573 4641 7607 4675
rect 7665 4641 7699 4675
rect 14841 4641 14875 4675
rect 5549 4573 5583 4607
rect 5733 4573 5767 4607
rect 6009 4573 6043 4607
rect 6193 4573 6227 4607
rect 7297 4573 7331 4607
rect 7481 4573 7515 4607
rect 7849 4573 7883 4607
rect 13277 4573 13311 4607
rect 13645 4573 13679 4607
rect 15025 4573 15059 4607
rect 15485 4573 15519 4607
rect 15669 4573 15703 4607
rect 15945 4573 15979 4607
rect 16405 4573 16439 4607
rect 16773 4573 16807 4607
rect 17049 4573 17083 4607
rect 18521 4573 18555 4607
rect 5365 4505 5399 4539
rect 17294 4505 17328 4539
rect 6101 4437 6135 4471
rect 8033 4437 8067 4471
rect 13461 4437 13495 4471
rect 15209 4437 15243 4471
rect 16957 4437 16991 4471
rect 18429 4437 18463 4471
rect 18705 4437 18739 4471
rect 15209 4233 15243 4267
rect 16681 4233 16715 4267
rect 17601 4233 17635 4267
rect 17785 4233 17819 4267
rect 10977 4165 11011 4199
rect 11193 4165 11227 4199
rect 15945 4165 15979 4199
rect 16145 4165 16179 4199
rect 16833 4165 16867 4199
rect 17049 4165 17083 4199
rect 19174 4165 19208 4199
rect 4629 4097 4663 4131
rect 5181 4097 5215 4131
rect 5365 4097 5399 4131
rect 5457 4097 5491 4131
rect 6377 4097 6411 4131
rect 7389 4097 7423 4131
rect 8125 4097 8159 4131
rect 8217 4097 8251 4131
rect 8401 4097 8435 4131
rect 9413 4097 9447 4131
rect 9597 4097 9631 4131
rect 9965 4097 9999 4131
rect 11529 4097 11563 4131
rect 12918 4097 12952 4131
rect 13277 4097 13311 4131
rect 13829 4097 13863 4131
rect 14013 4097 14047 4131
rect 15853 4097 15887 4131
rect 17693 4097 17727 4131
rect 19441 4097 19475 4131
rect 20646 4097 20680 4131
rect 20913 4097 20947 4131
rect 4813 4029 4847 4063
rect 4905 4029 4939 4063
rect 6101 4029 6135 4063
rect 6929 4029 6963 4063
rect 9505 4029 9539 4063
rect 9781 4029 9815 4063
rect 13185 4029 13219 4063
rect 14197 4029 14231 4063
rect 14289 4029 14323 4063
rect 14841 4029 14875 4063
rect 17969 4029 18003 4063
rect 5549 3961 5583 3995
rect 8033 3961 8067 3995
rect 11345 3961 11379 3995
rect 11713 3961 11747 3995
rect 16313 3961 16347 3995
rect 4445 3893 4479 3927
rect 4997 3893 5031 3927
rect 8401 3893 8435 3927
rect 10149 3893 10183 3927
rect 11161 3893 11195 3927
rect 11805 3893 11839 3927
rect 13461 3893 13495 3927
rect 16129 3893 16163 3927
rect 16865 3893 16899 3927
rect 17417 3893 17451 3927
rect 18061 3893 18095 3927
rect 19533 3893 19567 3927
rect 7205 3689 7239 3723
rect 7389 3689 7423 3723
rect 8677 3689 8711 3723
rect 9505 3689 9539 3723
rect 9965 3689 9999 3723
rect 12449 3689 12483 3723
rect 12909 3689 12943 3723
rect 13369 3689 13403 3723
rect 16313 3689 16347 3723
rect 16497 3689 16531 3723
rect 17417 3689 17451 3723
rect 17877 3689 17911 3723
rect 18705 3689 18739 3723
rect 20177 3689 20211 3723
rect 6377 3621 6411 3655
rect 7021 3621 7055 3655
rect 8585 3621 8619 3655
rect 10333 3621 10367 3655
rect 10517 3621 10551 3655
rect 10701 3621 10735 3655
rect 15485 3621 15519 3655
rect 17325 3621 17359 3655
rect 7113 3553 7147 3587
rect 8309 3553 8343 3587
rect 8769 3553 8803 3587
rect 12541 3553 12575 3587
rect 14105 3553 14139 3587
rect 16129 3553 16163 3587
rect 16957 3553 16991 3587
rect 18521 3553 18555 3587
rect 4997 3485 5031 3519
rect 6653 3485 6687 3519
rect 7665 3485 7699 3519
rect 8033 3485 8067 3519
rect 8125 3485 8159 3519
rect 8401 3485 8435 3519
rect 8493 3485 8527 3519
rect 9137 3485 9171 3519
rect 9597 3485 9631 3519
rect 9689 3485 9723 3519
rect 10057 3485 10091 3519
rect 10609 3485 10643 3519
rect 10793 3485 10827 3519
rect 11069 3485 11103 3519
rect 11621 3485 11655 3519
rect 11989 3485 12023 3519
rect 12081 3485 12115 3519
rect 12265 3485 12299 3519
rect 12357 3485 12391 3519
rect 12725 3485 12759 3519
rect 13001 3485 13035 3519
rect 13185 3485 13219 3519
rect 13645 3485 13679 3519
rect 13829 3485 13863 3519
rect 15577 3485 15611 3519
rect 16497 3485 16531 3519
rect 16589 3485 16623 3519
rect 16773 3485 16807 3519
rect 17141 3485 17175 3519
rect 17601 3485 17635 3519
rect 17693 3485 17727 3519
rect 17969 3485 18003 3519
rect 18889 3485 18923 3519
rect 19073 3485 19107 3519
rect 19257 3485 19291 3519
rect 19809 3485 19843 3519
rect 19993 3485 20027 3519
rect 5242 3417 5276 3451
rect 9321 3417 9355 3451
rect 11805 3417 11839 3451
rect 12449 3417 12483 3451
rect 14350 3417 14384 3451
rect 17877 3417 17911 3451
rect 7849 3349 7883 3383
rect 9781 3349 9815 3383
rect 10057 3349 10091 3383
rect 10885 3349 10919 3383
rect 13461 3349 13495 3383
rect 6009 3145 6043 3179
rect 6535 3145 6569 3179
rect 6837 3145 6871 3179
rect 8401 3145 8435 3179
rect 10333 3145 10367 3179
rect 11529 3145 11563 3179
rect 14289 3145 14323 3179
rect 16129 3145 16163 3179
rect 16681 3145 16715 3179
rect 20361 3145 20395 3179
rect 6745 3077 6779 3111
rect 7972 3077 8006 3111
rect 9220 3077 9254 3111
rect 12357 3077 12391 3111
rect 14924 3077 14958 3111
rect 4445 3009 4479 3043
rect 4701 3009 4735 3043
rect 5917 3009 5951 3043
rect 6101 3009 6135 3043
rect 8217 3009 8251 3043
rect 8309 3009 8343 3043
rect 8585 3009 8619 3043
rect 8953 3009 8987 3043
rect 10517 3009 10551 3043
rect 10609 3009 10643 3043
rect 11047 3009 11081 3043
rect 11345 3009 11379 3043
rect 11713 3009 11747 3043
rect 11897 3009 11931 3043
rect 11989 3009 12023 3043
rect 12173 3009 12207 3043
rect 12449 3009 12483 3043
rect 12909 3009 12943 3043
rect 13176 3009 13210 3043
rect 14657 3009 14691 3043
rect 16313 3009 16347 3043
rect 17794 3009 17828 3043
rect 18061 3009 18095 3043
rect 19266 3009 19300 3043
rect 19533 3009 19567 3043
rect 20177 3009 20211 3043
rect 11161 2941 11195 2975
rect 19993 2941 20027 2975
rect 5825 2873 5859 2907
rect 10977 2873 11011 2907
rect 11253 2873 11287 2907
rect 12173 2873 12207 2907
rect 16037 2873 16071 2907
rect 6377 2805 6411 2839
rect 6561 2805 6595 2839
rect 8585 2805 8619 2839
rect 18153 2805 18187 2839
rect 13369 2601 13403 2635
rect 17141 2601 17175 2635
rect 18889 2601 18923 2635
rect 19257 2601 19291 2635
rect 21465 2601 21499 2635
rect 18521 2465 18555 2499
rect 1409 2397 1443 2431
rect 9045 2397 9079 2431
rect 13553 2397 13587 2431
rect 16957 2397 16991 2431
rect 17417 2397 17451 2431
rect 17601 2397 17635 2431
rect 17785 2397 17819 2431
rect 17969 2397 18003 2431
rect 18705 2397 18739 2431
rect 19441 2397 19475 2431
rect 21649 2397 21683 2431
rect 1593 2261 1627 2295
rect 9137 2261 9171 2295
<< metal1 >>
rect 1104 22874 22264 22896
rect 1104 22822 4255 22874
rect 4307 22822 4319 22874
rect 4371 22822 4383 22874
rect 4435 22822 4447 22874
rect 4499 22822 4511 22874
rect 4563 22822 9545 22874
rect 9597 22822 9609 22874
rect 9661 22822 9673 22874
rect 9725 22822 9737 22874
rect 9789 22822 9801 22874
rect 9853 22822 14835 22874
rect 14887 22822 14899 22874
rect 14951 22822 14963 22874
rect 15015 22822 15027 22874
rect 15079 22822 15091 22874
rect 15143 22822 20125 22874
rect 20177 22822 20189 22874
rect 20241 22822 20253 22874
rect 20305 22822 20317 22874
rect 20369 22822 20381 22874
rect 20433 22822 22264 22874
rect 1104 22800 22264 22822
rect 1302 22720 1308 22772
rect 1360 22760 1366 22772
rect 1489 22763 1547 22769
rect 1489 22760 1501 22763
rect 1360 22732 1501 22760
rect 1360 22720 1366 22732
rect 1489 22729 1501 22732
rect 1535 22729 1547 22763
rect 1489 22723 1547 22729
rect 10318 22720 10324 22772
rect 10376 22760 10382 22772
rect 10689 22763 10747 22769
rect 10689 22760 10701 22763
rect 10376 22732 10701 22760
rect 10376 22720 10382 22732
rect 10689 22729 10701 22732
rect 10735 22729 10747 22763
rect 10689 22723 10747 22729
rect 19334 22720 19340 22772
rect 19392 22720 19398 22772
rect 1762 22584 1768 22636
rect 1820 22584 1826 22636
rect 10873 22627 10931 22633
rect 10873 22593 10885 22627
rect 10919 22624 10931 22627
rect 13265 22627 13323 22633
rect 13265 22624 13277 22627
rect 10919 22596 13277 22624
rect 10919 22593 10931 22596
rect 10873 22587 10931 22593
rect 13265 22593 13277 22596
rect 13311 22593 13323 22627
rect 13265 22587 13323 22593
rect 13446 22584 13452 22636
rect 13504 22584 13510 22636
rect 13630 22584 13636 22636
rect 13688 22584 13694 22636
rect 13725 22627 13783 22633
rect 13725 22593 13737 22627
rect 13771 22593 13783 22627
rect 13725 22587 13783 22593
rect 13538 22516 13544 22568
rect 13596 22556 13602 22568
rect 13740 22556 13768 22587
rect 16758 22584 16764 22636
rect 16816 22584 16822 22636
rect 19352 22624 19380 22720
rect 19613 22627 19671 22633
rect 19613 22624 19625 22627
rect 19352 22596 19625 22624
rect 19613 22593 19625 22596
rect 19659 22593 19671 22627
rect 19613 22587 19671 22593
rect 13596 22528 13768 22556
rect 13596 22516 13602 22528
rect 16942 22380 16948 22432
rect 17000 22380 17006 22432
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 19429 22423 19487 22429
rect 19429 22420 19441 22423
rect 19392 22392 19441 22420
rect 19392 22380 19398 22392
rect 19429 22389 19441 22392
rect 19475 22389 19487 22423
rect 19429 22383 19487 22389
rect 1104 22330 22264 22352
rect 1104 22278 3595 22330
rect 3647 22278 3659 22330
rect 3711 22278 3723 22330
rect 3775 22278 3787 22330
rect 3839 22278 3851 22330
rect 3903 22278 8885 22330
rect 8937 22278 8949 22330
rect 9001 22278 9013 22330
rect 9065 22278 9077 22330
rect 9129 22278 9141 22330
rect 9193 22278 14175 22330
rect 14227 22278 14239 22330
rect 14291 22278 14303 22330
rect 14355 22278 14367 22330
rect 14419 22278 14431 22330
rect 14483 22278 19465 22330
rect 19517 22278 19529 22330
rect 19581 22278 19593 22330
rect 19645 22278 19657 22330
rect 19709 22278 19721 22330
rect 19773 22278 22264 22330
rect 1104 22256 22264 22278
rect 7469 22219 7527 22225
rect 7469 22185 7481 22219
rect 7515 22216 7527 22219
rect 7515 22188 8432 22216
rect 7515 22185 7527 22188
rect 7469 22179 7527 22185
rect 8404 22160 8432 22188
rect 7377 22151 7435 22157
rect 7377 22117 7389 22151
rect 7423 22148 7435 22151
rect 7558 22148 7564 22160
rect 7423 22120 7564 22148
rect 7423 22117 7435 22120
rect 7377 22111 7435 22117
rect 7558 22108 7564 22120
rect 7616 22108 7622 22160
rect 8386 22108 8392 22160
rect 8444 22108 8450 22160
rect 12986 22108 12992 22160
rect 13044 22148 13050 22160
rect 13541 22151 13599 22157
rect 13541 22148 13553 22151
rect 13044 22120 13553 22148
rect 13044 22108 13050 22120
rect 13541 22117 13553 22120
rect 13587 22117 13599 22151
rect 13541 22111 13599 22117
rect 2590 22040 2596 22092
rect 2648 22080 2654 22092
rect 4890 22080 4896 22092
rect 2648 22052 4896 22080
rect 2648 22040 2654 22052
rect 4890 22040 4896 22052
rect 4948 22080 4954 22092
rect 5169 22083 5227 22089
rect 5169 22080 5181 22083
rect 4948 22052 5181 22080
rect 4948 22040 4954 22052
rect 5169 22049 5181 22052
rect 5215 22049 5227 22083
rect 7469 22083 7527 22089
rect 7469 22080 7481 22083
rect 5169 22043 5227 22049
rect 6748 22052 7481 22080
rect 6748 22024 6776 22052
rect 7469 22049 7481 22052
rect 7515 22049 7527 22083
rect 12710 22080 12716 22092
rect 7469 22043 7527 22049
rect 11992 22052 12716 22080
rect 3237 22015 3295 22021
rect 3237 21981 3249 22015
rect 3283 22012 3295 22015
rect 3418 22012 3424 22024
rect 3283 21984 3424 22012
rect 3283 21981 3295 21984
rect 3237 21975 3295 21981
rect 3418 21972 3424 21984
rect 3476 21972 3482 22024
rect 4341 22015 4399 22021
rect 4341 22012 4353 22015
rect 4080 21984 4353 22012
rect 2958 21904 2964 21956
rect 3016 21904 3022 21956
rect 4080 21888 4108 21984
rect 4341 21981 4353 21984
rect 4387 21981 4399 22015
rect 4341 21975 4399 21981
rect 6730 21972 6736 22024
rect 6788 21972 6794 22024
rect 7285 22015 7343 22021
rect 7285 21981 7297 22015
rect 7331 21981 7343 22015
rect 7285 21975 7343 21981
rect 7745 22015 7803 22021
rect 7745 21981 7757 22015
rect 7791 21981 7803 22015
rect 7745 21975 7803 21981
rect 5436 21947 5494 21953
rect 5436 21913 5448 21947
rect 5482 21944 5494 21947
rect 5718 21944 5724 21956
rect 5482 21916 5724 21944
rect 5482 21913 5494 21916
rect 5436 21907 5494 21913
rect 5718 21904 5724 21916
rect 5776 21904 5782 21956
rect 7300 21944 7328 21975
rect 7374 21944 7380 21956
rect 7300 21916 7380 21944
rect 7374 21904 7380 21916
rect 7432 21904 7438 21956
rect 7653 21947 7711 21953
rect 7653 21913 7665 21947
rect 7699 21913 7711 21947
rect 7653 21907 7711 21913
rect 3050 21836 3056 21888
rect 3108 21885 3114 21888
rect 3108 21839 3117 21885
rect 3145 21879 3203 21885
rect 3145 21845 3157 21879
rect 3191 21876 3203 21879
rect 3510 21876 3516 21888
rect 3191 21848 3516 21876
rect 3191 21845 3203 21848
rect 3145 21839 3203 21845
rect 3108 21836 3114 21839
rect 3510 21836 3516 21848
rect 3568 21876 3574 21888
rect 3789 21879 3847 21885
rect 3789 21876 3801 21879
rect 3568 21848 3801 21876
rect 3568 21836 3574 21848
rect 3789 21845 3801 21848
rect 3835 21845 3847 21879
rect 3789 21839 3847 21845
rect 4062 21836 4068 21888
rect 4120 21836 4126 21888
rect 6549 21879 6607 21885
rect 6549 21845 6561 21879
rect 6595 21876 6607 21879
rect 7098 21876 7104 21888
rect 6595 21848 7104 21876
rect 6595 21845 6607 21848
rect 6549 21839 6607 21845
rect 7098 21836 7104 21848
rect 7156 21836 7162 21888
rect 7190 21836 7196 21888
rect 7248 21876 7254 21888
rect 7668 21876 7696 21907
rect 7760 21888 7788 21975
rect 8294 21972 8300 22024
rect 8352 21972 8358 22024
rect 9950 21972 9956 22024
rect 10008 21972 10014 22024
rect 11992 22021 12020 22052
rect 12710 22040 12716 22052
rect 12768 22080 12774 22092
rect 13265 22083 13323 22089
rect 13265 22080 13277 22083
rect 12768 22052 13277 22080
rect 12768 22040 12774 22052
rect 13265 22049 13277 22052
rect 13311 22049 13323 22083
rect 13265 22043 13323 22049
rect 11977 22015 12035 22021
rect 11977 22012 11989 22015
rect 11348 21984 11989 22012
rect 10220 21947 10278 21953
rect 10220 21913 10232 21947
rect 10266 21944 10278 21947
rect 10410 21944 10416 21956
rect 10266 21916 10416 21944
rect 10266 21913 10278 21916
rect 10220 21907 10278 21913
rect 10410 21904 10416 21916
rect 10468 21904 10474 21956
rect 7248 21848 7696 21876
rect 7248 21836 7254 21848
rect 7742 21836 7748 21888
rect 7800 21836 7806 21888
rect 7834 21836 7840 21888
rect 7892 21836 7898 21888
rect 8478 21836 8484 21888
rect 8536 21836 8542 21888
rect 11348 21885 11376 21984
rect 11977 21981 11989 21984
rect 12023 21981 12035 22015
rect 11977 21975 12035 21981
rect 12066 21972 12072 22024
rect 12124 22012 12130 22024
rect 12437 22015 12495 22021
rect 12437 22012 12449 22015
rect 12124 21984 12449 22012
rect 12124 21972 12130 21984
rect 12437 21981 12449 21984
rect 12483 21981 12495 22015
rect 12437 21975 12495 21981
rect 13078 21972 13084 22024
rect 13136 21972 13142 22024
rect 13556 22012 13584 22111
rect 15473 22015 15531 22021
rect 13556 21984 15332 22012
rect 12158 21904 12164 21956
rect 12216 21904 12222 21956
rect 12342 21944 12348 21956
rect 12303 21916 12348 21944
rect 12342 21904 12348 21916
rect 12400 21944 12406 21956
rect 12529 21947 12587 21953
rect 12529 21944 12541 21947
rect 12400 21916 12541 21944
rect 12400 21904 12406 21916
rect 12529 21913 12541 21916
rect 12575 21913 12587 21947
rect 12529 21907 12587 21913
rect 13648 21916 14136 21944
rect 13648 21888 13676 21916
rect 11333 21879 11391 21885
rect 11333 21845 11345 21879
rect 11379 21845 11391 21879
rect 11333 21839 11391 21845
rect 11422 21836 11428 21888
rect 11480 21836 11486 21888
rect 12066 21836 12072 21888
rect 12124 21876 12130 21888
rect 12259 21879 12317 21885
rect 12259 21876 12271 21879
rect 12124 21848 12271 21876
rect 12124 21836 12130 21848
rect 12259 21845 12271 21848
rect 12305 21845 12317 21879
rect 12259 21839 12317 21845
rect 13630 21836 13636 21888
rect 13688 21836 13694 21888
rect 13722 21836 13728 21888
rect 13780 21836 13786 21888
rect 14108 21885 14136 21916
rect 14274 21904 14280 21956
rect 14332 21944 14338 21956
rect 15206 21947 15264 21953
rect 15206 21944 15218 21947
rect 14332 21916 15218 21944
rect 14332 21904 14338 21916
rect 15206 21913 15218 21916
rect 15252 21913 15264 21947
rect 15206 21907 15264 21913
rect 15304 21888 15332 21984
rect 15473 21981 15485 22015
rect 15519 22012 15531 22015
rect 17865 22015 17923 22021
rect 17865 22012 17877 22015
rect 15519 21984 17877 22012
rect 15519 21981 15531 21984
rect 15473 21975 15531 21981
rect 17865 21981 17877 21984
rect 17911 22012 17923 22015
rect 19058 22012 19064 22024
rect 17911 21984 19064 22012
rect 17911 21981 17923 21984
rect 17865 21975 17923 21981
rect 19058 21972 19064 21984
rect 19116 21972 19122 22024
rect 16942 21904 16948 21956
rect 17000 21944 17006 21956
rect 17598 21947 17656 21953
rect 17598 21944 17610 21947
rect 17000 21916 17610 21944
rect 17000 21904 17006 21916
rect 17598 21913 17610 21916
rect 17644 21913 17656 21947
rect 17598 21907 17656 21913
rect 14093 21879 14151 21885
rect 14093 21845 14105 21879
rect 14139 21845 14151 21879
rect 14093 21839 14151 21845
rect 15286 21836 15292 21888
rect 15344 21876 15350 21888
rect 16485 21879 16543 21885
rect 16485 21876 16497 21879
rect 15344 21848 16497 21876
rect 15344 21836 15350 21848
rect 16485 21845 16497 21848
rect 16531 21845 16543 21879
rect 16485 21839 16543 21845
rect 1104 21786 22264 21808
rect 1104 21734 4255 21786
rect 4307 21734 4319 21786
rect 4371 21734 4383 21786
rect 4435 21734 4447 21786
rect 4499 21734 4511 21786
rect 4563 21734 9545 21786
rect 9597 21734 9609 21786
rect 9661 21734 9673 21786
rect 9725 21734 9737 21786
rect 9789 21734 9801 21786
rect 9853 21734 14835 21786
rect 14887 21734 14899 21786
rect 14951 21734 14963 21786
rect 15015 21734 15027 21786
rect 15079 21734 15091 21786
rect 15143 21734 20125 21786
rect 20177 21734 20189 21786
rect 20241 21734 20253 21786
rect 20305 21734 20317 21786
rect 20369 21734 20381 21786
rect 20433 21734 22264 21786
rect 1104 21712 22264 21734
rect 2608 21644 2774 21672
rect 2317 21539 2375 21545
rect 2317 21505 2329 21539
rect 2363 21505 2375 21539
rect 2317 21499 2375 21505
rect 1762 21428 1768 21480
rect 1820 21428 1826 21480
rect 2332 21468 2360 21499
rect 2498 21496 2504 21548
rect 2556 21496 2562 21548
rect 2608 21545 2636 21644
rect 2593 21539 2651 21545
rect 2593 21505 2605 21539
rect 2639 21505 2651 21539
rect 2746 21536 2774 21644
rect 3050 21632 3056 21684
rect 3108 21632 3114 21684
rect 5718 21632 5724 21684
rect 5776 21632 5782 21684
rect 5997 21675 6055 21681
rect 5997 21641 6009 21675
rect 6043 21672 6055 21675
rect 6822 21672 6828 21684
rect 6043 21644 6828 21672
rect 6043 21641 6055 21644
rect 5997 21635 6055 21641
rect 6822 21632 6828 21644
rect 6880 21632 6886 21684
rect 6917 21675 6975 21681
rect 6917 21641 6929 21675
rect 6963 21672 6975 21675
rect 7190 21672 7196 21684
rect 6963 21644 7196 21672
rect 6963 21641 6975 21644
rect 6917 21635 6975 21641
rect 7190 21632 7196 21644
rect 7248 21632 7254 21684
rect 10410 21632 10416 21684
rect 10468 21632 10474 21684
rect 11422 21632 11428 21684
rect 11480 21632 11486 21684
rect 11882 21632 11888 21684
rect 11940 21632 11946 21684
rect 12066 21632 12072 21684
rect 12124 21632 12130 21684
rect 13078 21632 13084 21684
rect 13136 21632 13142 21684
rect 13173 21675 13231 21681
rect 13173 21641 13185 21675
rect 13219 21672 13231 21675
rect 13446 21672 13452 21684
rect 13219 21644 13452 21672
rect 13219 21641 13231 21644
rect 13173 21635 13231 21641
rect 13446 21632 13452 21644
rect 13504 21632 13510 21684
rect 13722 21632 13728 21684
rect 13780 21632 13786 21684
rect 14274 21632 14280 21684
rect 14332 21632 14338 21684
rect 15028 21644 16068 21672
rect 2952 21607 3010 21613
rect 2952 21573 2964 21607
rect 2998 21604 3010 21607
rect 3068 21604 3096 21632
rect 2998 21576 3096 21604
rect 5169 21607 5227 21613
rect 2998 21573 3010 21576
rect 2952 21567 3010 21573
rect 5169 21573 5181 21607
rect 5215 21604 5227 21607
rect 6086 21604 6092 21616
rect 5215 21576 6092 21604
rect 5215 21573 5227 21576
rect 5169 21567 5227 21573
rect 6086 21564 6092 21576
rect 6144 21564 6150 21616
rect 7834 21604 7840 21616
rect 6839 21576 7840 21604
rect 5353 21539 5411 21545
rect 2746 21508 4108 21536
rect 2593 21499 2651 21505
rect 2685 21471 2743 21477
rect 2332 21440 2544 21468
rect 1780 21400 1808 21428
rect 2317 21403 2375 21409
rect 2317 21400 2329 21403
rect 1780 21372 2329 21400
rect 2317 21369 2329 21372
rect 2363 21369 2375 21403
rect 2317 21363 2375 21369
rect 2516 21332 2544 21440
rect 2685 21437 2697 21471
rect 2731 21437 2743 21471
rect 2685 21431 2743 21437
rect 2590 21360 2596 21412
rect 2648 21400 2654 21412
rect 2700 21400 2728 21431
rect 4080 21412 4108 21508
rect 5353 21505 5365 21539
rect 5399 21505 5411 21539
rect 5353 21499 5411 21505
rect 5537 21539 5595 21545
rect 5537 21505 5549 21539
rect 5583 21536 5595 21539
rect 5721 21539 5779 21545
rect 5583 21508 5672 21536
rect 5583 21505 5595 21508
rect 5537 21499 5595 21505
rect 5368 21468 5396 21499
rect 5368 21440 5580 21468
rect 2648 21372 2728 21400
rect 2648 21360 2654 21372
rect 4062 21360 4068 21412
rect 4120 21360 4126 21412
rect 5552 21344 5580 21440
rect 5644 21400 5672 21508
rect 5721 21505 5733 21539
rect 5767 21505 5779 21539
rect 5721 21499 5779 21505
rect 5736 21468 5764 21499
rect 6178 21496 6184 21548
rect 6236 21496 6242 21548
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21536 6607 21539
rect 6730 21536 6736 21548
rect 6595 21508 6736 21536
rect 6595 21505 6607 21508
rect 6549 21499 6607 21505
rect 6730 21496 6736 21508
rect 6788 21496 6794 21548
rect 6839 21545 6867 21576
rect 7834 21564 7840 21576
rect 7892 21564 7898 21616
rect 8478 21564 8484 21616
rect 8536 21604 8542 21616
rect 9134 21607 9192 21613
rect 9134 21604 9146 21607
rect 8536 21576 9146 21604
rect 8536 21564 8542 21576
rect 9134 21573 9146 21576
rect 9180 21573 9192 21607
rect 11440 21604 11468 21632
rect 9134 21567 9192 21573
rect 10888 21576 11468 21604
rect 6825 21539 6883 21545
rect 6825 21505 6837 21539
rect 6871 21505 6883 21539
rect 6825 21499 6883 21505
rect 7098 21496 7104 21548
rect 7156 21536 7162 21548
rect 10888 21545 10916 21576
rect 7653 21539 7711 21545
rect 7653 21536 7665 21539
rect 7156 21508 7665 21536
rect 7156 21496 7162 21508
rect 7653 21505 7665 21508
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 10597 21539 10655 21545
rect 10597 21505 10609 21539
rect 10643 21505 10655 21539
rect 10597 21499 10655 21505
rect 10873 21539 10931 21545
rect 10873 21505 10885 21539
rect 10919 21505 10931 21539
rect 10873 21499 10931 21505
rect 6270 21468 6276 21480
rect 5736 21440 6276 21468
rect 6270 21428 6276 21440
rect 6328 21428 6334 21480
rect 6641 21471 6699 21477
rect 6641 21437 6653 21471
rect 6687 21468 6699 21471
rect 6914 21468 6920 21480
rect 6687 21440 6920 21468
rect 6687 21437 6699 21440
rect 6641 21431 6699 21437
rect 6914 21428 6920 21440
rect 6972 21468 6978 21480
rect 7558 21468 7564 21480
rect 6972 21440 7564 21468
rect 6972 21428 6978 21440
rect 7558 21428 7564 21440
rect 7616 21428 7622 21480
rect 9401 21471 9459 21477
rect 9401 21437 9413 21471
rect 9447 21468 9459 21471
rect 10612 21468 10640 21499
rect 10962 21496 10968 21548
rect 11020 21496 11026 21548
rect 11149 21539 11207 21545
rect 11149 21505 11161 21539
rect 11195 21536 11207 21539
rect 11900 21536 11928 21632
rect 11968 21607 12026 21613
rect 11968 21573 11980 21607
rect 12014 21604 12026 21607
rect 12084 21604 12112 21632
rect 13740 21604 13768 21632
rect 12014 21576 12112 21604
rect 13372 21576 13768 21604
rect 12014 21573 12026 21576
rect 11968 21567 12026 21573
rect 13372 21545 13400 21576
rect 11195 21508 11928 21536
rect 13357 21539 13415 21545
rect 11195 21505 11207 21508
rect 11149 21499 11207 21505
rect 13357 21505 13369 21539
rect 13403 21505 13415 21539
rect 13357 21499 13415 21505
rect 13446 21496 13452 21548
rect 13504 21496 13510 21548
rect 13630 21496 13636 21548
rect 13688 21536 13694 21548
rect 15028 21545 15056 21644
rect 15197 21607 15255 21613
rect 15197 21573 15209 21607
rect 15243 21604 15255 21607
rect 15286 21604 15292 21616
rect 15243 21576 15292 21604
rect 15243 21573 15255 21576
rect 15197 21567 15255 21573
rect 15286 21564 15292 21576
rect 15344 21564 15350 21616
rect 13725 21539 13783 21545
rect 13725 21536 13737 21539
rect 13688 21508 13737 21536
rect 13688 21496 13694 21508
rect 13725 21505 13737 21508
rect 13771 21536 13783 21539
rect 14553 21539 14611 21545
rect 14553 21536 14565 21539
rect 13771 21508 14565 21536
rect 13771 21505 13783 21508
rect 13725 21499 13783 21505
rect 14553 21505 14565 21508
rect 14599 21505 14611 21539
rect 15013 21539 15071 21545
rect 15013 21536 15025 21539
rect 14553 21499 14611 21505
rect 14660 21508 15025 21536
rect 11057 21471 11115 21477
rect 11057 21468 11069 21471
rect 9447 21440 9674 21468
rect 10612 21440 11069 21468
rect 9447 21437 9459 21440
rect 9401 21431 9459 21437
rect 5718 21400 5724 21412
rect 5644 21372 5724 21400
rect 5718 21360 5724 21372
rect 5776 21360 5782 21412
rect 8021 21403 8079 21409
rect 8021 21400 8033 21403
rect 6656 21372 8033 21400
rect 6656 21344 6684 21372
rect 8021 21369 8033 21372
rect 8067 21369 8079 21403
rect 8021 21363 8079 21369
rect 3970 21332 3976 21344
rect 2516 21304 3976 21332
rect 3970 21292 3976 21304
rect 4028 21292 4034 21344
rect 5534 21292 5540 21344
rect 5592 21292 5598 21344
rect 5813 21335 5871 21341
rect 5813 21301 5825 21335
rect 5859 21332 5871 21335
rect 6365 21335 6423 21341
rect 6365 21332 6377 21335
rect 5859 21304 6377 21332
rect 5859 21301 5871 21304
rect 5813 21295 5871 21301
rect 6365 21301 6377 21304
rect 6411 21301 6423 21335
rect 6365 21295 6423 21301
rect 6638 21292 6644 21344
rect 6696 21292 6702 21344
rect 6730 21292 6736 21344
rect 6788 21292 6794 21344
rect 7098 21292 7104 21344
rect 7156 21292 7162 21344
rect 9646 21332 9674 21440
rect 11057 21437 11069 21440
rect 11103 21437 11115 21471
rect 11057 21431 11115 21437
rect 11701 21471 11759 21477
rect 11701 21437 11713 21471
rect 11747 21437 11759 21471
rect 11701 21431 11759 21437
rect 11716 21400 11744 21431
rect 13538 21428 13544 21480
rect 13596 21428 13602 21480
rect 13909 21471 13967 21477
rect 13909 21437 13921 21471
rect 13955 21437 13967 21471
rect 13909 21431 13967 21437
rect 9876 21372 11744 21400
rect 13556 21400 13584 21428
rect 13633 21403 13691 21409
rect 13633 21400 13645 21403
rect 13556 21372 13645 21400
rect 9876 21344 9904 21372
rect 13633 21369 13645 21372
rect 13679 21369 13691 21403
rect 13924 21400 13952 21431
rect 13998 21428 14004 21480
rect 14056 21428 14062 21480
rect 14090 21428 14096 21480
rect 14148 21428 14154 21480
rect 14660 21477 14688 21508
rect 15013 21505 15025 21508
rect 15059 21505 15071 21539
rect 15304 21536 15332 21564
rect 16040 21548 16068 21644
rect 16574 21632 16580 21684
rect 16632 21672 16638 21684
rect 17129 21675 17187 21681
rect 16632 21644 17080 21672
rect 16632 21632 16638 21644
rect 17052 21604 17080 21644
rect 17129 21641 17141 21675
rect 17175 21672 17187 21675
rect 17379 21675 17437 21681
rect 17379 21672 17391 21675
rect 17175 21644 17391 21672
rect 17175 21641 17187 21644
rect 17129 21635 17187 21641
rect 17379 21641 17391 21644
rect 17425 21641 17437 21675
rect 17379 21635 17437 21641
rect 17589 21607 17647 21613
rect 17589 21604 17601 21607
rect 16316 21576 16988 21604
rect 17052 21576 17601 21604
rect 15838 21536 15844 21548
rect 15304 21508 15844 21536
rect 15013 21499 15071 21505
rect 14645 21471 14703 21477
rect 14645 21437 14657 21471
rect 14691 21437 14703 21471
rect 15028 21468 15056 21499
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 16022 21496 16028 21548
rect 16080 21496 16086 21548
rect 16114 21496 16120 21548
rect 16172 21496 16178 21548
rect 15194 21468 15200 21480
rect 15028 21440 15200 21468
rect 14645 21431 14703 21437
rect 15194 21428 15200 21440
rect 15252 21428 15258 21480
rect 15286 21428 15292 21480
rect 15344 21468 15350 21480
rect 16316 21477 16344 21576
rect 16485 21539 16543 21545
rect 16485 21505 16497 21539
rect 16531 21536 16543 21539
rect 16666 21536 16672 21548
rect 16531 21508 16672 21536
rect 16531 21505 16543 21508
rect 16485 21499 16543 21505
rect 16666 21496 16672 21508
rect 16724 21496 16730 21548
rect 16960 21545 16988 21576
rect 17589 21573 17601 21576
rect 17635 21573 17647 21607
rect 17589 21567 17647 21573
rect 16945 21539 17003 21545
rect 16945 21505 16957 21539
rect 16991 21505 17003 21539
rect 16945 21499 17003 21505
rect 21637 21539 21695 21545
rect 21637 21505 21649 21539
rect 21683 21536 21695 21539
rect 22186 21536 22192 21548
rect 21683 21508 22192 21536
rect 21683 21505 21695 21508
rect 21637 21499 21695 21505
rect 22186 21496 22192 21508
rect 22244 21496 22250 21548
rect 16301 21471 16359 21477
rect 16301 21468 16313 21471
rect 15344 21440 16313 21468
rect 15344 21428 15350 21440
rect 16301 21437 16313 21440
rect 16347 21437 16359 21471
rect 16761 21471 16819 21477
rect 16761 21468 16773 21471
rect 16301 21431 16359 21437
rect 16408 21440 16773 21468
rect 15010 21400 15016 21412
rect 13924 21372 15016 21400
rect 13633 21363 13691 21369
rect 15010 21360 15016 21372
rect 15068 21360 15074 21412
rect 16025 21403 16083 21409
rect 16025 21369 16037 21403
rect 16071 21400 16083 21403
rect 16209 21403 16267 21409
rect 16209 21400 16221 21403
rect 16071 21372 16221 21400
rect 16071 21369 16083 21372
rect 16025 21363 16083 21369
rect 16209 21369 16221 21372
rect 16255 21400 16267 21403
rect 16408 21400 16436 21440
rect 16761 21437 16773 21440
rect 16807 21437 16819 21471
rect 16761 21431 16819 21437
rect 16255 21372 16436 21400
rect 16255 21369 16267 21372
rect 16209 21363 16267 21369
rect 16942 21360 16948 21412
rect 17000 21400 17006 21412
rect 17000 21372 17448 21400
rect 17000 21360 17006 21372
rect 9858 21332 9864 21344
rect 9646 21304 9864 21332
rect 9858 21292 9864 21304
rect 9916 21292 9922 21344
rect 10778 21292 10784 21344
rect 10836 21292 10842 21344
rect 14918 21292 14924 21344
rect 14976 21292 14982 21344
rect 15381 21335 15439 21341
rect 15381 21301 15393 21335
rect 15427 21332 15439 21335
rect 15470 21332 15476 21344
rect 15427 21304 15476 21332
rect 15427 21301 15439 21304
rect 15381 21295 15439 21301
rect 15470 21292 15476 21304
rect 15528 21292 15534 21344
rect 16298 21292 16304 21344
rect 16356 21292 16362 21344
rect 16758 21292 16764 21344
rect 16816 21292 16822 21344
rect 16850 21292 16856 21344
rect 16908 21332 16914 21344
rect 17420 21341 17448 21372
rect 17221 21335 17279 21341
rect 17221 21332 17233 21335
rect 16908 21304 17233 21332
rect 16908 21292 16914 21304
rect 17221 21301 17233 21304
rect 17267 21301 17279 21335
rect 17221 21295 17279 21301
rect 17405 21335 17463 21341
rect 17405 21301 17417 21335
rect 17451 21301 17463 21335
rect 17405 21295 17463 21301
rect 20622 21292 20628 21344
rect 20680 21332 20686 21344
rect 21453 21335 21511 21341
rect 21453 21332 21465 21335
rect 20680 21304 21465 21332
rect 20680 21292 20686 21304
rect 21453 21301 21465 21304
rect 21499 21301 21511 21335
rect 21453 21295 21511 21301
rect 1104 21242 22264 21264
rect 1104 21190 3595 21242
rect 3647 21190 3659 21242
rect 3711 21190 3723 21242
rect 3775 21190 3787 21242
rect 3839 21190 3851 21242
rect 3903 21190 8885 21242
rect 8937 21190 8949 21242
rect 9001 21190 9013 21242
rect 9065 21190 9077 21242
rect 9129 21190 9141 21242
rect 9193 21190 14175 21242
rect 14227 21190 14239 21242
rect 14291 21190 14303 21242
rect 14355 21190 14367 21242
rect 14419 21190 14431 21242
rect 14483 21190 19465 21242
rect 19517 21190 19529 21242
rect 19581 21190 19593 21242
rect 19645 21190 19657 21242
rect 19709 21190 19721 21242
rect 19773 21190 22264 21242
rect 1104 21168 22264 21190
rect 2498 21088 2504 21140
rect 2556 21088 2562 21140
rect 2958 21088 2964 21140
rect 3016 21128 3022 21140
rect 3329 21131 3387 21137
rect 3329 21128 3341 21131
rect 3016 21100 3341 21128
rect 3016 21088 3022 21100
rect 3329 21097 3341 21100
rect 3375 21097 3387 21131
rect 3329 21091 3387 21097
rect 3418 21088 3424 21140
rect 3476 21088 3482 21140
rect 3510 21088 3516 21140
rect 3568 21088 3574 21140
rect 3789 21131 3847 21137
rect 3789 21097 3801 21131
rect 3835 21128 3847 21131
rect 3970 21128 3976 21140
rect 3835 21100 3976 21128
rect 3835 21097 3847 21100
rect 3789 21091 3847 21097
rect 3970 21088 3976 21100
rect 4028 21088 4034 21140
rect 4062 21088 4068 21140
rect 4120 21128 4126 21140
rect 4249 21131 4307 21137
rect 4249 21128 4261 21131
rect 4120 21100 4261 21128
rect 4120 21088 4126 21100
rect 4249 21097 4261 21100
rect 4295 21097 4307 21131
rect 4249 21091 4307 21097
rect 6178 21088 6184 21140
rect 6236 21088 6242 21140
rect 6270 21088 6276 21140
rect 6328 21088 6334 21140
rect 6365 21131 6423 21137
rect 6365 21097 6377 21131
rect 6411 21128 6423 21131
rect 6730 21128 6736 21140
rect 6411 21100 6736 21128
rect 6411 21097 6423 21100
rect 6365 21091 6423 21097
rect 6730 21088 6736 21100
rect 6788 21088 6794 21140
rect 6822 21088 6828 21140
rect 6880 21088 6886 21140
rect 7009 21131 7067 21137
rect 7009 21097 7021 21131
rect 7055 21128 7067 21131
rect 7374 21128 7380 21140
rect 7055 21100 7380 21128
rect 7055 21097 7067 21100
rect 7009 21091 7067 21097
rect 7374 21088 7380 21100
rect 7432 21128 7438 21140
rect 7742 21128 7748 21140
rect 7432 21100 7748 21128
rect 7432 21088 7438 21100
rect 7742 21088 7748 21100
rect 7800 21088 7806 21140
rect 7834 21088 7840 21140
rect 7892 21088 7898 21140
rect 8294 21088 8300 21140
rect 8352 21088 8358 21140
rect 8478 21088 8484 21140
rect 8536 21088 8542 21140
rect 9677 21131 9735 21137
rect 9677 21097 9689 21131
rect 9723 21128 9735 21131
rect 10410 21128 10416 21140
rect 9723 21100 10416 21128
rect 9723 21097 9735 21100
rect 9677 21091 9735 21097
rect 10410 21088 10416 21100
rect 10468 21088 10474 21140
rect 11974 21088 11980 21140
rect 12032 21088 12038 21140
rect 12161 21131 12219 21137
rect 12161 21097 12173 21131
rect 12207 21128 12219 21131
rect 12250 21128 12256 21140
rect 12207 21100 12256 21128
rect 12207 21097 12219 21100
rect 12161 21091 12219 21097
rect 2516 20856 2544 21088
rect 3237 20995 3295 21001
rect 3237 20961 3249 20995
rect 3283 20961 3295 20995
rect 3237 20955 3295 20961
rect 3142 20884 3148 20936
rect 3200 20924 3206 20936
rect 3252 20924 3280 20955
rect 3528 20933 3556 21088
rect 5813 21063 5871 21069
rect 5813 21029 5825 21063
rect 5859 21060 5871 21063
rect 6196 21060 6224 21088
rect 5859 21032 6224 21060
rect 6288 21060 6316 21088
rect 6840 21060 6868 21088
rect 7101 21063 7159 21069
rect 7101 21060 7113 21063
rect 6288 21032 6776 21060
rect 6840 21032 7113 21060
rect 5859 21029 5871 21032
rect 5813 21023 5871 21029
rect 5534 20992 5540 21004
rect 4356 20964 5540 20992
rect 3200 20896 3280 20924
rect 3513 20927 3571 20933
rect 3200 20884 3206 20896
rect 3513 20893 3525 20927
rect 3559 20893 3571 20927
rect 3513 20887 3571 20893
rect 3970 20884 3976 20936
rect 4028 20884 4034 20936
rect 4062 20884 4068 20936
rect 4120 20884 4126 20936
rect 4356 20933 4384 20964
rect 5534 20952 5540 20964
rect 5592 20992 5598 21004
rect 5997 20995 6055 21001
rect 5592 20964 5948 20992
rect 5592 20952 5598 20964
rect 5920 20936 5948 20964
rect 5997 20961 6009 20995
rect 6043 20992 6055 20995
rect 6086 20992 6092 21004
rect 6043 20964 6092 20992
rect 6043 20961 6055 20964
rect 5997 20955 6055 20961
rect 6086 20952 6092 20964
rect 6144 20952 6150 21004
rect 4341 20927 4399 20933
rect 4341 20893 4353 20927
rect 4387 20893 4399 20927
rect 4341 20887 4399 20893
rect 5721 20927 5779 20933
rect 5721 20893 5733 20927
rect 5767 20924 5779 20927
rect 5810 20924 5816 20936
rect 5767 20896 5816 20924
rect 5767 20893 5779 20896
rect 5721 20887 5779 20893
rect 4356 20856 4384 20887
rect 5810 20884 5816 20896
rect 5868 20884 5874 20936
rect 5902 20884 5908 20936
rect 5960 20884 5966 20936
rect 6196 20933 6224 21032
rect 6638 20952 6644 21004
rect 6696 20952 6702 21004
rect 6748 20992 6776 21032
rect 7101 21029 7113 21032
rect 7147 21029 7159 21063
rect 7852 21060 7880 21088
rect 7101 21023 7159 21029
rect 7484 21032 7880 21060
rect 11149 21063 11207 21069
rect 6748 20964 7236 20992
rect 6181 20927 6239 20933
rect 6181 20893 6193 20927
rect 6227 20893 6239 20927
rect 6181 20887 6239 20893
rect 6825 20927 6883 20933
rect 6825 20893 6837 20927
rect 6871 20893 6883 20927
rect 6825 20887 6883 20893
rect 2516 20828 4384 20856
rect 6840 20800 6868 20887
rect 5810 20748 5816 20800
rect 5868 20788 5874 20800
rect 6822 20788 6828 20800
rect 5868 20760 6828 20788
rect 5868 20748 5874 20760
rect 6822 20748 6828 20760
rect 6880 20748 6886 20800
rect 7208 20788 7236 20964
rect 7484 20933 7512 21032
rect 11149 21029 11161 21063
rect 11195 21060 11207 21063
rect 11195 21032 11928 21060
rect 11195 21029 11207 21032
rect 11149 21023 11207 21029
rect 11900 21001 11928 21032
rect 7837 20995 7895 21001
rect 7837 20992 7849 20995
rect 7576 20964 7849 20992
rect 7576 20936 7604 20964
rect 7837 20961 7849 20964
rect 7883 20961 7895 20995
rect 7837 20955 7895 20961
rect 11885 20995 11943 21001
rect 11885 20961 11897 20995
rect 11931 20992 11943 20995
rect 12176 20992 12204 21091
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 12710 21088 12716 21140
rect 12768 21088 12774 21140
rect 12986 21088 12992 21140
rect 13044 21088 13050 21140
rect 13078 21088 13084 21140
rect 13136 21088 13142 21140
rect 13357 21131 13415 21137
rect 13357 21097 13369 21131
rect 13403 21128 13415 21131
rect 13538 21128 13544 21140
rect 13403 21100 13544 21128
rect 13403 21097 13415 21100
rect 13357 21091 13415 21097
rect 13538 21088 13544 21100
rect 13596 21088 13602 21140
rect 14090 21088 14096 21140
rect 14148 21128 14154 21140
rect 14737 21131 14795 21137
rect 14737 21128 14749 21131
rect 14148 21100 14749 21128
rect 14148 21088 14154 21100
rect 14737 21097 14749 21100
rect 14783 21097 14795 21131
rect 14737 21091 14795 21097
rect 14918 21088 14924 21140
rect 14976 21088 14982 21140
rect 15010 21088 15016 21140
rect 15068 21128 15074 21140
rect 15381 21131 15439 21137
rect 15381 21128 15393 21131
rect 15068 21100 15393 21128
rect 15068 21088 15074 21100
rect 15381 21097 15393 21100
rect 15427 21097 15439 21131
rect 15381 21091 15439 21097
rect 15470 21088 15476 21140
rect 15528 21128 15534 21140
rect 15528 21100 15700 21128
rect 15528 21088 15534 21100
rect 11931 20964 12204 20992
rect 11931 20961 11943 20964
rect 11885 20955 11943 20961
rect 7450 20927 7512 20933
rect 7299 20905 7357 20911
rect 7299 20871 7311 20905
rect 7345 20902 7357 20905
rect 7345 20874 7420 20902
rect 7450 20893 7462 20927
rect 7496 20896 7512 20927
rect 7496 20893 7508 20896
rect 7450 20887 7508 20893
rect 7558 20884 7564 20936
rect 7616 20884 7622 20936
rect 7650 20884 7656 20936
rect 7708 20924 7714 20936
rect 8021 20927 8079 20933
rect 8021 20924 8033 20927
rect 7708 20896 8033 20924
rect 7708 20884 7714 20896
rect 8021 20893 8033 20896
rect 8067 20893 8079 20927
rect 8021 20887 8079 20893
rect 9493 20927 9551 20933
rect 9493 20893 9505 20927
rect 9539 20893 9551 20927
rect 9493 20887 9551 20893
rect 9677 20927 9735 20933
rect 9677 20893 9689 20927
rect 9723 20893 9735 20927
rect 9677 20887 9735 20893
rect 9769 20927 9827 20933
rect 9769 20893 9781 20927
rect 9815 20924 9827 20927
rect 9858 20924 9864 20936
rect 9815 20896 9864 20924
rect 9815 20893 9827 20896
rect 9769 20887 9827 20893
rect 7345 20871 7357 20874
rect 7299 20865 7357 20871
rect 7392 20856 7420 20874
rect 7742 20856 7748 20868
rect 7392 20828 7748 20856
rect 7742 20816 7748 20828
rect 7800 20816 7806 20868
rect 8128 20828 8616 20856
rect 8128 20788 8156 20828
rect 7208 20760 8156 20788
rect 8205 20791 8263 20797
rect 8205 20757 8217 20791
rect 8251 20788 8263 20791
rect 8455 20791 8513 20797
rect 8455 20788 8467 20791
rect 8251 20760 8467 20788
rect 8251 20757 8263 20760
rect 8205 20751 8263 20757
rect 8455 20757 8467 20760
rect 8501 20757 8513 20791
rect 8588 20788 8616 20828
rect 8662 20816 8668 20868
rect 8720 20816 8726 20868
rect 9306 20788 9312 20800
rect 8588 20760 9312 20788
rect 8455 20751 8513 20757
rect 9306 20748 9312 20760
rect 9364 20748 9370 20800
rect 9508 20788 9536 20887
rect 9692 20856 9720 20887
rect 9858 20884 9864 20896
rect 9916 20884 9922 20936
rect 10778 20924 10784 20936
rect 9968 20896 10784 20924
rect 9968 20856 9996 20896
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 12728 20933 12756 21088
rect 12713 20927 12771 20933
rect 12713 20924 12725 20927
rect 12360 20896 12725 20924
rect 9692 20828 9996 20856
rect 10036 20859 10094 20865
rect 10036 20825 10048 20859
rect 10082 20856 10094 20859
rect 10226 20856 10232 20868
rect 10082 20828 10232 20856
rect 10082 20825 10094 20828
rect 10036 20819 10094 20825
rect 10226 20816 10232 20828
rect 10284 20816 10290 20868
rect 12360 20865 12388 20896
rect 12713 20893 12725 20896
rect 12759 20893 12771 20927
rect 13096 20924 13124 21088
rect 14936 20933 14964 21088
rect 15562 21060 15568 21072
rect 15028 21032 15568 21060
rect 15028 20933 15056 21032
rect 15562 21020 15568 21032
rect 15620 21020 15626 21072
rect 15672 21001 15700 21100
rect 15838 21088 15844 21140
rect 15896 21088 15902 21140
rect 16114 21088 16120 21140
rect 16172 21128 16178 21140
rect 16390 21128 16396 21140
rect 16172 21100 16396 21128
rect 16172 21088 16178 21100
rect 16390 21088 16396 21100
rect 16448 21128 16454 21140
rect 16758 21128 16764 21140
rect 16448 21100 16764 21128
rect 16448 21088 16454 21100
rect 16758 21088 16764 21100
rect 16816 21128 16822 21140
rect 17037 21131 17095 21137
rect 17037 21128 17049 21131
rect 16816 21100 17049 21128
rect 16816 21088 16822 21100
rect 17037 21097 17049 21100
rect 17083 21097 17095 21131
rect 17037 21091 17095 21097
rect 15657 20995 15715 21001
rect 15657 20992 15669 20995
rect 15120 20964 15669 20992
rect 15120 20933 15148 20964
rect 15657 20961 15669 20964
rect 15703 20961 15715 20995
rect 15657 20955 15715 20961
rect 15746 20952 15752 21004
rect 15804 20952 15810 21004
rect 15856 20992 15884 21088
rect 16022 21020 16028 21072
rect 16080 21060 16086 21072
rect 16080 21032 16896 21060
rect 16080 21020 16086 21032
rect 16669 20995 16727 21001
rect 16669 20992 16681 20995
rect 15856 20964 16681 20992
rect 16669 20961 16681 20964
rect 16715 20961 16727 20995
rect 16669 20955 16727 20961
rect 13265 20927 13323 20933
rect 13265 20924 13277 20927
rect 13096 20896 13277 20924
rect 12713 20887 12771 20893
rect 13265 20893 13277 20896
rect 13311 20893 13323 20927
rect 13265 20887 13323 20893
rect 14921 20927 14979 20933
rect 14921 20893 14933 20927
rect 14967 20893 14979 20927
rect 14921 20887 14979 20893
rect 15013 20927 15071 20933
rect 15013 20893 15025 20927
rect 15059 20893 15071 20927
rect 15013 20887 15071 20893
rect 15105 20927 15163 20933
rect 15105 20893 15117 20927
rect 15151 20893 15163 20927
rect 15105 20887 15163 20893
rect 15212 20896 15516 20924
rect 12129 20859 12187 20865
rect 12129 20856 12141 20859
rect 11164 20828 12141 20856
rect 11164 20800 11192 20828
rect 12129 20825 12141 20828
rect 12175 20825 12187 20859
rect 12129 20819 12187 20825
rect 12345 20859 12403 20865
rect 12345 20825 12357 20859
rect 12391 20825 12403 20859
rect 14936 20856 14964 20887
rect 15212 20856 15240 20896
rect 14936 20828 15240 20856
rect 15289 20859 15347 20865
rect 12345 20819 12403 20825
rect 15289 20825 15301 20859
rect 15335 20825 15347 20859
rect 15488 20856 15516 20896
rect 15562 20884 15568 20936
rect 15620 20884 15626 20936
rect 16868 20933 16896 21032
rect 15841 20927 15899 20933
rect 15841 20893 15853 20927
rect 15887 20893 15899 20927
rect 15841 20887 15899 20893
rect 16853 20927 16911 20933
rect 16853 20893 16865 20927
rect 16899 20893 16911 20927
rect 16853 20887 16911 20893
rect 15856 20856 15884 20887
rect 15488 20828 15884 20856
rect 15289 20819 15347 20825
rect 10318 20788 10324 20800
rect 9508 20760 10324 20788
rect 10318 20748 10324 20760
rect 10376 20788 10382 20800
rect 10962 20788 10968 20800
rect 10376 20760 10968 20788
rect 10376 20748 10382 20760
rect 10962 20748 10968 20760
rect 11020 20748 11026 20800
rect 11146 20748 11152 20800
rect 11204 20748 11210 20800
rect 11238 20748 11244 20800
rect 11296 20748 11302 20800
rect 13078 20748 13084 20800
rect 13136 20788 13142 20800
rect 13173 20791 13231 20797
rect 13173 20788 13185 20791
rect 13136 20760 13185 20788
rect 13136 20748 13142 20760
rect 13173 20757 13185 20760
rect 13219 20757 13231 20791
rect 15304 20788 15332 20819
rect 15470 20788 15476 20800
rect 15304 20760 15476 20788
rect 13173 20751 13231 20757
rect 15470 20748 15476 20760
rect 15528 20788 15534 20800
rect 15746 20788 15752 20800
rect 15528 20760 15752 20788
rect 15528 20748 15534 20760
rect 15746 20748 15752 20760
rect 15804 20748 15810 20800
rect 1104 20698 22264 20720
rect 1104 20646 4255 20698
rect 4307 20646 4319 20698
rect 4371 20646 4383 20698
rect 4435 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 9545 20698
rect 9597 20646 9609 20698
rect 9661 20646 9673 20698
rect 9725 20646 9737 20698
rect 9789 20646 9801 20698
rect 9853 20646 14835 20698
rect 14887 20646 14899 20698
rect 14951 20646 14963 20698
rect 15015 20646 15027 20698
rect 15079 20646 15091 20698
rect 15143 20646 20125 20698
rect 20177 20646 20189 20698
rect 20241 20646 20253 20698
rect 20305 20646 20317 20698
rect 20369 20646 20381 20698
rect 20433 20646 22264 20698
rect 1104 20624 22264 20646
rect 3881 20587 3939 20593
rect 3881 20553 3893 20587
rect 3927 20584 3939 20587
rect 3970 20584 3976 20596
rect 3927 20556 3976 20584
rect 3927 20553 3939 20556
rect 3881 20547 3939 20553
rect 3970 20544 3976 20556
rect 4028 20544 4034 20596
rect 5902 20544 5908 20596
rect 5960 20584 5966 20596
rect 6549 20587 6607 20593
rect 6549 20584 6561 20587
rect 5960 20556 6561 20584
rect 5960 20544 5966 20556
rect 6549 20553 6561 20556
rect 6595 20553 6607 20587
rect 6549 20547 6607 20553
rect 6825 20587 6883 20593
rect 6825 20553 6837 20587
rect 6871 20584 6883 20587
rect 6914 20584 6920 20596
rect 6871 20556 6920 20584
rect 6871 20553 6883 20556
rect 6825 20547 6883 20553
rect 6914 20544 6920 20556
rect 6972 20544 6978 20596
rect 7098 20544 7104 20596
rect 7156 20544 7162 20596
rect 7282 20544 7288 20596
rect 7340 20584 7346 20596
rect 7742 20584 7748 20596
rect 7340 20556 7748 20584
rect 7340 20544 7346 20556
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 10226 20544 10232 20596
rect 10284 20544 10290 20596
rect 10778 20544 10784 20596
rect 10836 20544 10842 20596
rect 11977 20587 12035 20593
rect 11977 20553 11989 20587
rect 12023 20584 12035 20587
rect 12158 20584 12164 20596
rect 12023 20556 12164 20584
rect 12023 20553 12035 20556
rect 11977 20547 12035 20553
rect 12158 20544 12164 20556
rect 12216 20544 12222 20596
rect 12250 20544 12256 20596
rect 12308 20584 12314 20596
rect 12308 20556 12434 20584
rect 12308 20544 12314 20556
rect 7116 20516 7144 20544
rect 6656 20488 7144 20516
rect 6656 20457 6684 20488
rect 8662 20476 8668 20528
rect 8720 20516 8726 20528
rect 9033 20519 9091 20525
rect 9033 20516 9045 20519
rect 8720 20488 9045 20516
rect 8720 20476 8726 20488
rect 9033 20485 9045 20488
rect 9079 20516 9091 20519
rect 11330 20516 11336 20528
rect 9079 20488 11336 20516
rect 9079 20485 9091 20488
rect 9033 20479 9091 20485
rect 11330 20476 11336 20488
rect 11388 20476 11394 20528
rect 12406 20516 12434 20556
rect 15286 20544 15292 20596
rect 15344 20544 15350 20596
rect 15562 20544 15568 20596
rect 15620 20584 15626 20596
rect 15841 20587 15899 20593
rect 15841 20584 15853 20587
rect 15620 20556 15853 20584
rect 15620 20544 15626 20556
rect 15841 20553 15853 20556
rect 15887 20553 15899 20587
rect 15841 20547 15899 20553
rect 16040 20556 16988 20584
rect 11716 20488 12480 20516
rect 6641 20451 6699 20457
rect 6641 20417 6653 20451
rect 6687 20417 6699 20451
rect 6641 20411 6699 20417
rect 6730 20408 6736 20460
rect 6788 20408 6794 20460
rect 6822 20408 6828 20460
rect 6880 20448 6886 20460
rect 6917 20451 6975 20457
rect 6917 20448 6929 20451
rect 6880 20420 6929 20448
rect 6880 20408 6886 20420
rect 6917 20417 6929 20420
rect 6963 20417 6975 20451
rect 6917 20411 6975 20417
rect 10410 20408 10416 20460
rect 10468 20408 10474 20460
rect 10962 20408 10968 20460
rect 11020 20408 11026 20460
rect 11238 20448 11244 20460
rect 11072 20420 11244 20448
rect 3421 20383 3479 20389
rect 3421 20349 3433 20383
rect 3467 20380 3479 20383
rect 6748 20380 6776 20408
rect 3467 20352 6776 20380
rect 10689 20383 10747 20389
rect 3467 20349 3479 20352
rect 3421 20343 3479 20349
rect 10689 20349 10701 20383
rect 10735 20380 10747 20383
rect 11072 20380 11100 20420
rect 11238 20408 11244 20420
rect 11296 20408 11302 20460
rect 10735 20352 11100 20380
rect 11149 20383 11207 20389
rect 10735 20349 10747 20352
rect 10689 20343 10747 20349
rect 11149 20349 11161 20383
rect 11195 20380 11207 20383
rect 11716 20380 11744 20488
rect 12066 20408 12072 20460
rect 12124 20448 12130 20460
rect 12161 20451 12219 20457
rect 12161 20448 12173 20451
rect 12124 20420 12173 20448
rect 12124 20408 12130 20420
rect 12161 20417 12173 20420
rect 12207 20417 12219 20451
rect 12161 20411 12219 20417
rect 12253 20451 12311 20457
rect 12253 20417 12265 20451
rect 12299 20448 12311 20451
rect 12342 20448 12348 20460
rect 12299 20420 12348 20448
rect 12299 20417 12311 20420
rect 12253 20411 12311 20417
rect 12342 20408 12348 20420
rect 12400 20408 12406 20460
rect 12452 20457 12480 20488
rect 12437 20451 12495 20457
rect 12437 20417 12449 20451
rect 12483 20417 12495 20451
rect 12437 20411 12495 20417
rect 15194 20408 15200 20460
rect 15252 20408 15258 20460
rect 15378 20408 15384 20460
rect 15436 20408 15442 20460
rect 15746 20408 15752 20460
rect 15804 20408 15810 20460
rect 16040 20457 16068 20556
rect 16132 20488 16896 20516
rect 16132 20460 16160 20488
rect 16025 20451 16083 20457
rect 16025 20417 16037 20451
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 16114 20408 16120 20460
rect 16172 20408 16178 20460
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20417 16359 20451
rect 16301 20411 16359 20417
rect 11195 20352 11744 20380
rect 11977 20383 12035 20389
rect 11195 20349 11207 20352
rect 11149 20343 11207 20349
rect 11977 20349 11989 20383
rect 12023 20380 12035 20383
rect 16206 20380 16212 20392
rect 12023 20352 16212 20380
rect 12023 20349 12035 20352
rect 11977 20343 12035 20349
rect 3789 20315 3847 20321
rect 3789 20281 3801 20315
rect 3835 20312 3847 20315
rect 3970 20312 3976 20324
rect 3835 20284 3976 20312
rect 3835 20281 3847 20284
rect 3789 20275 3847 20281
rect 3970 20272 3976 20284
rect 4028 20272 4034 20324
rect 11992 20312 12020 20343
rect 12268 20324 12296 20352
rect 16206 20340 16212 20352
rect 16264 20340 16270 20392
rect 16316 20380 16344 20411
rect 16390 20408 16396 20460
rect 16448 20408 16454 20460
rect 16868 20457 16896 20488
rect 16960 20460 16988 20556
rect 20622 20544 20628 20596
rect 20680 20544 20686 20596
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 16684 20380 16712 20411
rect 16942 20408 16948 20460
rect 17000 20408 17006 20460
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20448 20407 20451
rect 20640 20448 20668 20544
rect 20395 20420 20668 20448
rect 20395 20417 20407 20420
rect 20349 20411 20407 20417
rect 16316 20352 16712 20380
rect 20165 20383 20223 20389
rect 9140 20284 12020 20312
rect 3142 20204 3148 20256
rect 3200 20244 3206 20256
rect 9140 20253 9168 20284
rect 12250 20272 12256 20324
rect 12308 20272 12314 20324
rect 16408 20256 16436 20352
rect 20165 20349 20177 20383
rect 20211 20349 20223 20383
rect 20165 20343 20223 20349
rect 16666 20272 16672 20324
rect 16724 20272 16730 20324
rect 20180 20256 20208 20343
rect 9125 20247 9183 20253
rect 9125 20244 9137 20247
rect 3200 20216 9137 20244
rect 3200 20204 3206 20216
rect 9125 20213 9137 20216
rect 9171 20213 9183 20247
rect 9125 20207 9183 20213
rect 10597 20247 10655 20253
rect 10597 20213 10609 20247
rect 10643 20244 10655 20247
rect 11146 20244 11152 20256
rect 10643 20216 11152 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 11146 20204 11152 20216
rect 11204 20204 11210 20256
rect 12526 20204 12532 20256
rect 12584 20204 12590 20256
rect 15470 20204 15476 20256
rect 15528 20244 15534 20256
rect 15565 20247 15623 20253
rect 15565 20244 15577 20247
rect 15528 20216 15577 20244
rect 15528 20204 15534 20216
rect 15565 20213 15577 20216
rect 15611 20244 15623 20247
rect 16114 20244 16120 20256
rect 15611 20216 16120 20244
rect 15611 20213 15623 20216
rect 15565 20207 15623 20213
rect 16114 20204 16120 20216
rect 16172 20204 16178 20256
rect 16390 20204 16396 20256
rect 16448 20204 16454 20256
rect 20162 20204 20168 20256
rect 20220 20204 20226 20256
rect 20530 20204 20536 20256
rect 20588 20204 20594 20256
rect 1104 20154 22264 20176
rect 1104 20102 3595 20154
rect 3647 20102 3659 20154
rect 3711 20102 3723 20154
rect 3775 20102 3787 20154
rect 3839 20102 3851 20154
rect 3903 20102 8885 20154
rect 8937 20102 8949 20154
rect 9001 20102 9013 20154
rect 9065 20102 9077 20154
rect 9129 20102 9141 20154
rect 9193 20102 14175 20154
rect 14227 20102 14239 20154
rect 14291 20102 14303 20154
rect 14355 20102 14367 20154
rect 14419 20102 14431 20154
rect 14483 20102 19465 20154
rect 19517 20102 19529 20154
rect 19581 20102 19593 20154
rect 19645 20102 19657 20154
rect 19709 20102 19721 20154
rect 19773 20102 22264 20154
rect 1104 20080 22264 20102
rect 4709 20043 4767 20049
rect 4709 20040 4721 20043
rect 4356 20012 4721 20040
rect 2884 19876 3556 19904
rect 2884 19845 2912 19876
rect 3160 19845 3188 19876
rect 3528 19848 3556 19876
rect 2869 19839 2927 19845
rect 2869 19805 2881 19839
rect 2915 19805 2927 19839
rect 2869 19799 2927 19805
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19805 3111 19839
rect 3053 19799 3111 19805
rect 3145 19839 3203 19845
rect 3145 19805 3157 19839
rect 3191 19805 3203 19839
rect 3145 19799 3203 19805
rect 3068 19768 3096 19799
rect 3234 19796 3240 19848
rect 3292 19796 3298 19848
rect 3329 19839 3387 19845
rect 3329 19805 3341 19839
rect 3375 19836 3387 19839
rect 3418 19836 3424 19848
rect 3375 19808 3424 19836
rect 3375 19805 3387 19808
rect 3329 19799 3387 19805
rect 3418 19796 3424 19808
rect 3476 19796 3482 19848
rect 3510 19796 3516 19848
rect 3568 19796 3574 19848
rect 3970 19796 3976 19848
rect 4028 19836 4034 19848
rect 4356 19845 4384 20012
rect 4709 20009 4721 20012
rect 4755 20009 4767 20043
rect 4709 20003 4767 20009
rect 12526 20000 12532 20052
rect 12584 20000 12590 20052
rect 13446 20000 13452 20052
rect 13504 20040 13510 20052
rect 13725 20043 13783 20049
rect 13725 20040 13737 20043
rect 13504 20012 13737 20040
rect 13504 20000 13510 20012
rect 13725 20009 13737 20012
rect 13771 20009 13783 20043
rect 13725 20003 13783 20009
rect 15746 20000 15752 20052
rect 15804 20000 15810 20052
rect 16206 20000 16212 20052
rect 16264 20000 16270 20052
rect 16390 20000 16396 20052
rect 16448 20000 16454 20052
rect 16761 20043 16819 20049
rect 16761 20009 16773 20043
rect 16807 20040 16819 20043
rect 17402 20040 17408 20052
rect 16807 20012 17408 20040
rect 16807 20009 16819 20012
rect 16761 20003 16819 20009
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 20530 20000 20536 20052
rect 20588 20000 20594 20052
rect 12544 19904 12572 20000
rect 16224 19972 16252 20000
rect 20162 19972 20168 19984
rect 16224 19944 20168 19972
rect 13354 19904 13360 19916
rect 12544 19876 13360 19904
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 19628 19913 19656 19944
rect 20162 19932 20168 19944
rect 20220 19932 20226 19984
rect 16853 19907 16911 19913
rect 16853 19904 16865 19907
rect 13556 19876 16865 19904
rect 4341 19839 4399 19845
rect 4341 19836 4353 19839
rect 4028 19808 4353 19836
rect 4028 19796 4034 19808
rect 4341 19805 4353 19808
rect 4387 19805 4399 19839
rect 4341 19799 4399 19805
rect 4985 19839 5043 19845
rect 4985 19805 4997 19839
rect 5031 19836 5043 19839
rect 6730 19836 6736 19848
rect 5031 19808 6736 19836
rect 5031 19805 5043 19808
rect 4985 19799 5043 19805
rect 6730 19796 6736 19808
rect 6788 19796 6794 19848
rect 12894 19796 12900 19848
rect 12952 19796 12958 19848
rect 12989 19839 13047 19845
rect 12989 19805 13001 19839
rect 13035 19836 13047 19839
rect 13078 19836 13084 19848
rect 13035 19808 13084 19836
rect 13035 19805 13047 19808
rect 12989 19799 13047 19805
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13170 19796 13176 19848
rect 13228 19796 13234 19848
rect 13262 19796 13268 19848
rect 13320 19796 13326 19848
rect 13556 19845 13584 19876
rect 16853 19873 16865 19876
rect 16899 19873 16911 19907
rect 16853 19867 16911 19873
rect 17681 19907 17739 19913
rect 17681 19873 17693 19907
rect 17727 19873 17739 19907
rect 17681 19867 17739 19873
rect 19613 19907 19671 19913
rect 19613 19873 19625 19907
rect 19659 19873 19671 19907
rect 19613 19867 19671 19873
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 3252 19768 3280 19796
rect 12912 19768 12940 19796
rect 13556 19768 13584 19799
rect 15194 19796 15200 19848
rect 15252 19836 15258 19848
rect 15565 19839 15623 19845
rect 15565 19836 15577 19839
rect 15252 19808 15577 19836
rect 15252 19796 15258 19808
rect 15565 19805 15577 19808
rect 15611 19836 15623 19839
rect 16298 19836 16304 19848
rect 15611 19808 16304 19836
rect 15611 19805 15623 19808
rect 15565 19799 15623 19805
rect 16298 19796 16304 19808
rect 16356 19836 16362 19848
rect 16577 19839 16635 19845
rect 16577 19836 16589 19839
rect 16356 19808 16589 19836
rect 16356 19796 16362 19808
rect 16577 19805 16589 19808
rect 16623 19805 16635 19839
rect 16868 19836 16896 19867
rect 17586 19836 17592 19848
rect 16868 19808 17592 19836
rect 16577 19799 16635 19805
rect 3068 19740 4844 19768
rect 12912 19740 13584 19768
rect 4816 19712 4844 19740
rect 15378 19728 15384 19780
rect 15436 19728 15442 19780
rect 16592 19768 16620 19799
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 17696 19768 17724 19867
rect 19426 19796 19432 19848
rect 19484 19796 19490 19848
rect 20441 19839 20499 19845
rect 20441 19805 20453 19839
rect 20487 19836 20499 19839
rect 20548 19836 20576 20000
rect 20487 19808 20576 19836
rect 20487 19805 20499 19808
rect 20441 19799 20499 19805
rect 16592 19740 17724 19768
rect 2958 19660 2964 19712
rect 3016 19660 3022 19712
rect 3050 19660 3056 19712
rect 3108 19700 3114 19712
rect 3237 19703 3295 19709
rect 3237 19700 3249 19703
rect 3108 19672 3249 19700
rect 3108 19660 3114 19672
rect 3237 19669 3249 19672
rect 3283 19669 3295 19703
rect 3237 19663 3295 19669
rect 3418 19660 3424 19712
rect 3476 19700 3482 19712
rect 3789 19703 3847 19709
rect 3789 19700 3801 19703
rect 3476 19672 3801 19700
rect 3476 19660 3482 19672
rect 3789 19669 3801 19672
rect 3835 19669 3847 19703
rect 3789 19663 3847 19669
rect 4525 19703 4583 19709
rect 4525 19669 4537 19703
rect 4571 19700 4583 19703
rect 4614 19700 4620 19712
rect 4571 19672 4620 19700
rect 4571 19669 4583 19672
rect 4525 19663 4583 19669
rect 4614 19660 4620 19672
rect 4672 19660 4678 19712
rect 4798 19660 4804 19712
rect 4856 19660 4862 19712
rect 16022 19660 16028 19712
rect 16080 19700 16086 19712
rect 16758 19700 16764 19712
rect 16080 19672 16764 19700
rect 16080 19660 16086 19672
rect 16758 19660 16764 19672
rect 16816 19660 16822 19712
rect 17957 19703 18015 19709
rect 17957 19669 17969 19703
rect 18003 19700 18015 19703
rect 18138 19700 18144 19712
rect 18003 19672 18144 19700
rect 18003 19669 18015 19672
rect 17957 19663 18015 19669
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 19242 19660 19248 19712
rect 19300 19660 19306 19712
rect 20257 19703 20315 19709
rect 20257 19669 20269 19703
rect 20303 19700 20315 19703
rect 20622 19700 20628 19712
rect 20303 19672 20628 19700
rect 20303 19669 20315 19672
rect 20257 19663 20315 19669
rect 20622 19660 20628 19672
rect 20680 19660 20686 19712
rect 1104 19610 22264 19632
rect 1104 19558 4255 19610
rect 4307 19558 4319 19610
rect 4371 19558 4383 19610
rect 4435 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 9545 19610
rect 9597 19558 9609 19610
rect 9661 19558 9673 19610
rect 9725 19558 9737 19610
rect 9789 19558 9801 19610
rect 9853 19558 14835 19610
rect 14887 19558 14899 19610
rect 14951 19558 14963 19610
rect 15015 19558 15027 19610
rect 15079 19558 15091 19610
rect 15143 19558 20125 19610
rect 20177 19558 20189 19610
rect 20241 19558 20253 19610
rect 20305 19558 20317 19610
rect 20369 19558 20381 19610
rect 20433 19558 22264 19610
rect 1104 19536 22264 19558
rect 2777 19499 2835 19505
rect 2777 19465 2789 19499
rect 2823 19465 2835 19499
rect 2777 19459 2835 19465
rect 2590 19428 2596 19440
rect 1412 19400 2596 19428
rect 1412 19369 1440 19400
rect 2590 19388 2596 19400
rect 2648 19388 2654 19440
rect 2792 19428 2820 19459
rect 3326 19456 3332 19508
rect 3384 19496 3390 19508
rect 3421 19499 3479 19505
rect 3421 19496 3433 19499
rect 3384 19468 3433 19496
rect 3384 19456 3390 19468
rect 3421 19465 3433 19468
rect 3467 19465 3479 19499
rect 3970 19496 3976 19508
rect 3421 19459 3479 19465
rect 3528 19468 3976 19496
rect 3528 19428 3556 19468
rect 3804 19437 3832 19468
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 6822 19456 6828 19508
rect 6880 19496 6886 19508
rect 8570 19496 8576 19508
rect 6880 19468 8576 19496
rect 6880 19456 6886 19468
rect 8570 19456 8576 19468
rect 8628 19456 8634 19508
rect 12894 19456 12900 19508
rect 12952 19496 12958 19508
rect 12952 19468 13216 19496
rect 12952 19456 12958 19468
rect 2792 19400 3556 19428
rect 3589 19431 3647 19437
rect 3589 19397 3601 19431
rect 3635 19428 3647 19431
rect 3789 19431 3847 19437
rect 3635 19397 3648 19428
rect 3589 19391 3648 19397
rect 3789 19397 3801 19431
rect 3835 19397 3847 19431
rect 3789 19391 3847 19397
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19329 1455 19363
rect 1397 19323 1455 19329
rect 1664 19363 1722 19369
rect 1664 19329 1676 19363
rect 1710 19360 1722 19363
rect 2869 19363 2927 19369
rect 2869 19360 2881 19363
rect 1710 19332 2881 19360
rect 1710 19329 1722 19332
rect 1664 19323 1722 19329
rect 2869 19329 2881 19332
rect 2915 19329 2927 19363
rect 2869 19323 2927 19329
rect 3050 19320 3056 19372
rect 3108 19320 3114 19372
rect 3234 19320 3240 19372
rect 3292 19320 3298 19372
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 3418 19360 3424 19372
rect 3375 19332 3424 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 3418 19320 3424 19332
rect 3476 19320 3482 19372
rect 3252 19165 3280 19320
rect 3620 19224 3648 19391
rect 5994 19388 6000 19440
rect 6052 19428 6058 19440
rect 12713 19431 12771 19437
rect 6052 19400 7328 19428
rect 6052 19388 6058 19400
rect 5902 19320 5908 19372
rect 5960 19320 5966 19372
rect 6178 19320 6184 19372
rect 6236 19320 6242 19372
rect 6549 19363 6607 19369
rect 6549 19329 6561 19363
rect 6595 19360 6607 19363
rect 6822 19360 6828 19372
rect 6595 19332 6828 19360
rect 6595 19329 6607 19332
rect 6549 19323 6607 19329
rect 6822 19320 6828 19332
rect 6880 19320 6886 19372
rect 7300 19369 7328 19400
rect 10520 19400 11192 19428
rect 7009 19363 7067 19369
rect 7009 19329 7021 19363
rect 7055 19329 7067 19363
rect 7009 19323 7067 19329
rect 7285 19363 7343 19369
rect 7285 19329 7297 19363
rect 7331 19329 7343 19363
rect 7285 19323 7343 19329
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19360 7527 19363
rect 8113 19363 8171 19369
rect 7515 19332 8064 19360
rect 7515 19329 7527 19332
rect 7469 19323 7527 19329
rect 3344 19196 3648 19224
rect 6196 19224 6224 19320
rect 6270 19252 6276 19304
rect 6328 19292 6334 19304
rect 6365 19295 6423 19301
rect 6365 19292 6377 19295
rect 6328 19264 6377 19292
rect 6328 19252 6334 19264
rect 6365 19261 6377 19264
rect 6411 19292 6423 19295
rect 7024 19292 7052 19323
rect 6411 19264 7052 19292
rect 8036 19292 8064 19332
rect 8113 19329 8125 19363
rect 8159 19360 8171 19363
rect 9214 19360 9220 19372
rect 8159 19332 9220 19360
rect 8159 19329 8171 19332
rect 8113 19323 8171 19329
rect 9214 19320 9220 19332
rect 9272 19320 9278 19372
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19360 10379 19363
rect 10410 19360 10416 19372
rect 10367 19332 10416 19360
rect 10367 19329 10379 19332
rect 10321 19323 10379 19329
rect 10410 19320 10416 19332
rect 10468 19320 10474 19372
rect 10520 19369 10548 19400
rect 11164 19372 11192 19400
rect 12713 19397 12725 19431
rect 12759 19428 12771 19431
rect 12986 19428 12992 19440
rect 12759 19400 12992 19428
rect 12759 19397 12771 19400
rect 12713 19391 12771 19397
rect 12986 19388 12992 19400
rect 13044 19428 13050 19440
rect 13188 19437 13216 19468
rect 13262 19456 13268 19508
rect 13320 19496 13326 19508
rect 13449 19499 13507 19505
rect 13449 19496 13461 19499
rect 13320 19468 13461 19496
rect 13320 19456 13326 19468
rect 13449 19465 13461 19468
rect 13495 19465 13507 19499
rect 13449 19459 13507 19465
rect 16298 19456 16304 19508
rect 16356 19496 16362 19508
rect 16356 19468 16896 19496
rect 16356 19456 16362 19468
rect 13081 19431 13139 19437
rect 13081 19428 13093 19431
rect 13044 19400 13093 19428
rect 13044 19388 13050 19400
rect 13081 19397 13093 19400
rect 13127 19397 13139 19431
rect 13081 19391 13139 19397
rect 13173 19431 13231 19437
rect 13173 19397 13185 19431
rect 13219 19397 13231 19431
rect 13173 19391 13231 19397
rect 13354 19388 13360 19440
rect 13412 19388 13418 19440
rect 16868 19428 16896 19468
rect 17586 19456 17592 19508
rect 17644 19496 17650 19508
rect 17681 19499 17739 19505
rect 17681 19496 17693 19499
rect 17644 19468 17693 19496
rect 17644 19456 17650 19468
rect 17681 19465 17693 19468
rect 17727 19465 17739 19499
rect 17681 19459 17739 19465
rect 19242 19456 19248 19508
rect 19300 19456 19306 19508
rect 16868 19400 17632 19428
rect 10505 19363 10563 19369
rect 10505 19329 10517 19363
rect 10551 19329 10563 19363
rect 10505 19323 10563 19329
rect 11057 19363 11115 19369
rect 11057 19329 11069 19363
rect 11103 19329 11115 19363
rect 11057 19323 11115 19329
rect 8386 19292 8392 19304
rect 8036 19264 8392 19292
rect 6411 19261 6423 19264
rect 6365 19255 6423 19261
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 8662 19224 8668 19236
rect 6196 19196 8668 19224
rect 3344 19168 3372 19196
rect 8662 19184 8668 19196
rect 8720 19184 8726 19236
rect 11072 19224 11100 19323
rect 11146 19320 11152 19372
rect 11204 19320 11210 19372
rect 11882 19320 11888 19372
rect 11940 19320 11946 19372
rect 12618 19320 12624 19372
rect 12676 19320 12682 19372
rect 12897 19363 12955 19369
rect 12897 19329 12909 19363
rect 12943 19329 12955 19363
rect 12897 19323 12955 19329
rect 13265 19363 13323 19369
rect 13265 19329 13277 19363
rect 13311 19360 13323 19363
rect 13372 19360 13400 19388
rect 16657 19385 16715 19391
rect 16657 19382 16669 19385
rect 13311 19332 13400 19360
rect 13311 19329 13323 19332
rect 13265 19323 13323 19329
rect 11241 19295 11299 19301
rect 11241 19261 11253 19295
rect 11287 19292 11299 19295
rect 11974 19292 11980 19304
rect 11287 19264 11980 19292
rect 11287 19261 11299 19264
rect 11241 19255 11299 19261
rect 11974 19252 11980 19264
rect 12032 19292 12038 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 12032 19264 12449 19292
rect 12032 19252 12038 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12912 19292 12940 19323
rect 13538 19320 13544 19372
rect 13596 19320 13602 19372
rect 16298 19320 16304 19372
rect 16356 19320 16362 19372
rect 16485 19363 16543 19369
rect 16485 19329 16497 19363
rect 16531 19360 16543 19363
rect 16592 19360 16669 19382
rect 16531 19354 16669 19360
rect 16531 19332 16620 19354
rect 16657 19351 16669 19354
rect 16703 19351 16715 19385
rect 16657 19345 16715 19351
rect 16531 19329 16543 19332
rect 16485 19323 16543 19329
rect 16758 19320 16764 19372
rect 16816 19320 16822 19372
rect 17402 19360 17408 19372
rect 16868 19332 17408 19360
rect 13556 19292 13584 19320
rect 12912 19264 13584 19292
rect 16117 19295 16175 19301
rect 12437 19255 12495 19261
rect 16117 19261 16129 19295
rect 16163 19292 16175 19295
rect 16574 19292 16580 19304
rect 16163 19264 16580 19292
rect 16163 19261 16175 19264
rect 16117 19255 16175 19261
rect 16574 19252 16580 19264
rect 16632 19292 16638 19304
rect 16868 19292 16896 19332
rect 17402 19320 17408 19332
rect 17460 19320 17466 19372
rect 17604 19369 17632 19400
rect 17589 19363 17647 19369
rect 17589 19329 17601 19363
rect 17635 19329 17647 19363
rect 17589 19323 17647 19329
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 18794 19363 18852 19369
rect 18794 19360 18806 19363
rect 18380 19332 18806 19360
rect 18380 19320 18386 19332
rect 18794 19329 18806 19332
rect 18840 19329 18852 19363
rect 18794 19323 18852 19329
rect 19058 19320 19064 19372
rect 19116 19320 19122 19372
rect 19153 19363 19211 19369
rect 19153 19329 19165 19363
rect 19199 19360 19211 19363
rect 19260 19360 19288 19456
rect 19199 19332 19288 19360
rect 19199 19329 19211 19332
rect 19153 19323 19211 19329
rect 16632 19264 16896 19292
rect 16945 19295 17003 19301
rect 16632 19252 16638 19264
rect 16945 19261 16957 19295
rect 16991 19261 17003 19295
rect 16945 19255 17003 19261
rect 16960 19224 16988 19255
rect 17034 19252 17040 19304
rect 17092 19252 17098 19304
rect 19076 19292 19104 19320
rect 19334 19292 19340 19304
rect 19076 19264 19340 19292
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 17221 19227 17279 19233
rect 17221 19224 17233 19227
rect 11072 19196 12112 19224
rect 16960 19196 17233 19224
rect 12084 19168 12112 19196
rect 17221 19193 17233 19196
rect 17267 19193 17279 19227
rect 17221 19187 17279 19193
rect 3237 19159 3295 19165
rect 3237 19125 3249 19159
rect 3283 19125 3295 19159
rect 3237 19119 3295 19125
rect 3326 19116 3332 19168
rect 3384 19116 3390 19168
rect 3605 19159 3663 19165
rect 3605 19125 3617 19159
rect 3651 19156 3663 19159
rect 3970 19156 3976 19168
rect 3651 19128 3976 19156
rect 3651 19125 3663 19128
rect 3605 19119 3663 19125
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 6181 19159 6239 19165
rect 6181 19125 6193 19159
rect 6227 19156 6239 19159
rect 6546 19156 6552 19168
rect 6227 19128 6552 19156
rect 6227 19125 6239 19128
rect 6181 19119 6239 19125
rect 6546 19116 6552 19128
rect 6604 19116 6610 19168
rect 6638 19116 6644 19168
rect 6696 19156 6702 19168
rect 6733 19159 6791 19165
rect 6733 19156 6745 19159
rect 6696 19128 6745 19156
rect 6696 19116 6702 19128
rect 6733 19125 6745 19128
rect 6779 19125 6791 19159
rect 6733 19119 6791 19125
rect 7190 19116 7196 19168
rect 7248 19116 7254 19168
rect 7466 19116 7472 19168
rect 7524 19116 7530 19168
rect 7926 19116 7932 19168
rect 7984 19116 7990 19168
rect 8294 19116 8300 19168
rect 8352 19116 8358 19168
rect 10226 19116 10232 19168
rect 10284 19156 10290 19168
rect 10505 19159 10563 19165
rect 10505 19156 10517 19159
rect 10284 19128 10517 19156
rect 10284 19116 10290 19128
rect 10505 19125 10517 19128
rect 10551 19125 10563 19159
rect 10505 19119 10563 19125
rect 10870 19116 10876 19168
rect 10928 19116 10934 19168
rect 12066 19116 12072 19168
rect 12124 19116 12130 19168
rect 16206 19116 16212 19168
rect 16264 19156 16270 19168
rect 17034 19156 17040 19168
rect 16264 19128 17040 19156
rect 16264 19116 16270 19128
rect 17034 19116 17040 19128
rect 17092 19116 17098 19168
rect 17126 19116 17132 19168
rect 17184 19116 17190 19168
rect 19337 19159 19395 19165
rect 19337 19125 19349 19159
rect 19383 19156 19395 19159
rect 19886 19156 19892 19168
rect 19383 19128 19892 19156
rect 19383 19125 19395 19128
rect 19337 19119 19395 19125
rect 19886 19116 19892 19128
rect 19944 19116 19950 19168
rect 1104 19066 22264 19088
rect 1104 19014 3595 19066
rect 3647 19014 3659 19066
rect 3711 19014 3723 19066
rect 3775 19014 3787 19066
rect 3839 19014 3851 19066
rect 3903 19014 8885 19066
rect 8937 19014 8949 19066
rect 9001 19014 9013 19066
rect 9065 19014 9077 19066
rect 9129 19014 9141 19066
rect 9193 19014 14175 19066
rect 14227 19014 14239 19066
rect 14291 19014 14303 19066
rect 14355 19014 14367 19066
rect 14419 19014 14431 19066
rect 14483 19014 19465 19066
rect 19517 19014 19529 19066
rect 19581 19014 19593 19066
rect 19645 19014 19657 19066
rect 19709 19014 19721 19066
rect 19773 19014 22264 19066
rect 1104 18992 22264 19014
rect 2590 18952 2596 18964
rect 2240 18924 2596 18952
rect 2240 18825 2268 18924
rect 2590 18912 2596 18924
rect 2648 18912 2654 18964
rect 3789 18955 3847 18961
rect 3789 18921 3801 18955
rect 3835 18952 3847 18955
rect 4062 18952 4068 18964
rect 3835 18924 4068 18952
rect 3835 18921 3847 18924
rect 3789 18915 3847 18921
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 7650 18952 7656 18964
rect 7300 18924 7656 18952
rect 7300 18893 7328 18924
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 9214 18912 9220 18964
rect 9272 18912 9278 18964
rect 10321 18955 10379 18961
rect 10321 18921 10333 18955
rect 10367 18952 10379 18955
rect 10870 18952 10876 18964
rect 10367 18924 10876 18952
rect 10367 18921 10379 18924
rect 10321 18915 10379 18921
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 11885 18955 11943 18961
rect 11885 18921 11897 18955
rect 11931 18952 11943 18955
rect 11974 18952 11980 18964
rect 11931 18924 11980 18952
rect 11931 18921 11943 18924
rect 11885 18915 11943 18921
rect 11974 18912 11980 18924
rect 12032 18952 12038 18964
rect 12161 18955 12219 18961
rect 12161 18952 12173 18955
rect 12032 18924 12173 18952
rect 12032 18912 12038 18924
rect 12161 18921 12173 18924
rect 12207 18921 12219 18955
rect 12161 18915 12219 18921
rect 16025 18955 16083 18961
rect 16025 18921 16037 18955
rect 16071 18952 16083 18955
rect 16298 18952 16304 18964
rect 16071 18924 16304 18952
rect 16071 18921 16083 18924
rect 16025 18915 16083 18921
rect 16298 18912 16304 18924
rect 16356 18912 16362 18964
rect 16853 18955 16911 18961
rect 16853 18921 16865 18955
rect 16899 18952 16911 18955
rect 16942 18952 16948 18964
rect 16899 18924 16948 18952
rect 16899 18921 16911 18924
rect 16853 18915 16911 18921
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 17126 18912 17132 18964
rect 17184 18952 17190 18964
rect 17497 18955 17555 18961
rect 17497 18952 17509 18955
rect 17184 18924 17509 18952
rect 17184 18912 17190 18924
rect 17497 18921 17509 18924
rect 17543 18952 17555 18955
rect 17770 18952 17776 18964
rect 17543 18924 17776 18952
rect 17543 18921 17555 18924
rect 17497 18915 17555 18921
rect 17770 18912 17776 18924
rect 17828 18912 17834 18964
rect 17865 18955 17923 18961
rect 17865 18921 17877 18955
rect 17911 18952 17923 18955
rect 18322 18952 18328 18964
rect 17911 18924 18328 18952
rect 17911 18921 17923 18924
rect 17865 18915 17923 18921
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 7285 18887 7343 18893
rect 7285 18884 7297 18887
rect 6104 18856 7297 18884
rect 6104 18828 6132 18856
rect 7285 18853 7297 18856
rect 7331 18853 7343 18887
rect 16574 18884 16580 18896
rect 7285 18847 7343 18853
rect 15396 18856 16580 18884
rect 2225 18819 2283 18825
rect 2225 18785 2237 18819
rect 2271 18785 2283 18819
rect 4706 18816 4712 18828
rect 2225 18779 2283 18785
rect 3988 18788 4712 18816
rect 3988 18757 4016 18788
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 4890 18776 4896 18828
rect 4948 18776 4954 18828
rect 6086 18776 6092 18828
rect 6144 18776 6150 18828
rect 6656 18788 7052 18816
rect 3973 18751 4031 18757
rect 3973 18717 3985 18751
rect 4019 18717 4031 18751
rect 3973 18711 4031 18717
rect 4157 18751 4215 18757
rect 4157 18717 4169 18751
rect 4203 18717 4215 18751
rect 4157 18711 4215 18717
rect 4249 18751 4307 18757
rect 4249 18717 4261 18751
rect 4295 18717 4307 18751
rect 4249 18711 4307 18717
rect 4341 18751 4399 18757
rect 4341 18717 4353 18751
rect 4387 18717 4399 18751
rect 4341 18711 4399 18717
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18748 4583 18751
rect 4614 18748 4620 18760
rect 4571 18720 4620 18748
rect 4571 18717 4583 18720
rect 4525 18711 4583 18717
rect 2492 18683 2550 18689
rect 2492 18649 2504 18683
rect 2538 18680 2550 18683
rect 2774 18680 2780 18692
rect 2538 18652 2780 18680
rect 2538 18649 2550 18652
rect 2492 18643 2550 18649
rect 2774 18640 2780 18652
rect 2832 18640 2838 18692
rect 4172 18680 4200 18711
rect 3988 18652 4200 18680
rect 3988 18624 4016 18652
rect 3605 18615 3663 18621
rect 3605 18581 3617 18615
rect 3651 18612 3663 18615
rect 3970 18612 3976 18624
rect 3651 18584 3976 18612
rect 3651 18581 3663 18584
rect 3605 18575 3663 18581
rect 3970 18572 3976 18584
rect 4028 18572 4034 18624
rect 4154 18572 4160 18624
rect 4212 18612 4218 18624
rect 4264 18612 4292 18711
rect 4212 18584 4292 18612
rect 4356 18612 4384 18711
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18748 4859 18751
rect 6656 18748 6684 18788
rect 4847 18720 6684 18748
rect 4847 18717 4859 18720
rect 4801 18711 4859 18717
rect 6730 18708 6736 18760
rect 6788 18708 6794 18760
rect 5160 18683 5218 18689
rect 5160 18649 5172 18683
rect 5206 18680 5218 18683
rect 6362 18680 6368 18692
rect 5206 18652 6368 18680
rect 5206 18649 5218 18652
rect 5160 18643 5218 18649
rect 6362 18640 6368 18652
rect 6420 18640 6426 18692
rect 6457 18683 6515 18689
rect 6457 18649 6469 18683
rect 6503 18680 6515 18683
rect 6638 18680 6644 18692
rect 6503 18652 6644 18680
rect 6503 18649 6515 18652
rect 6457 18643 6515 18649
rect 6638 18640 6644 18652
rect 6696 18640 6702 18692
rect 4614 18612 4620 18624
rect 4356 18584 4620 18612
rect 4212 18572 4218 18584
rect 4614 18572 4620 18584
rect 4672 18572 4678 18624
rect 5534 18572 5540 18624
rect 5592 18612 5598 18624
rect 6270 18612 6276 18624
rect 5592 18584 6276 18612
rect 5592 18572 5598 18584
rect 6270 18572 6276 18584
rect 6328 18572 6334 18624
rect 7024 18612 7052 18788
rect 7190 18776 7196 18828
rect 7248 18776 7254 18828
rect 8386 18776 8392 18828
rect 8444 18816 8450 18828
rect 8846 18816 8852 18828
rect 8444 18788 8852 18816
rect 8444 18776 8450 18788
rect 8846 18776 8852 18788
rect 8904 18816 8910 18828
rect 10505 18819 10563 18825
rect 10505 18816 10517 18819
rect 8904 18788 9076 18816
rect 8904 18776 8910 18788
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 7208 18748 7236 18776
rect 7147 18720 7236 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 7374 18708 7380 18760
rect 7432 18708 7438 18760
rect 7644 18751 7702 18757
rect 7644 18717 7656 18751
rect 7690 18748 7702 18751
rect 7926 18748 7932 18760
rect 7690 18720 7932 18748
rect 7690 18717 7702 18720
rect 7644 18711 7702 18717
rect 7926 18708 7932 18720
rect 7984 18708 7990 18760
rect 9048 18757 9076 18788
rect 9968 18788 10517 18816
rect 9968 18760 9996 18788
rect 10505 18785 10517 18788
rect 10551 18785 10563 18819
rect 10505 18779 10563 18785
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8312 18720 8953 18748
rect 8312 18692 8340 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9033 18751 9091 18757
rect 9033 18717 9045 18751
rect 9079 18717 9091 18751
rect 9033 18711 9091 18717
rect 9950 18708 9956 18760
rect 10008 18708 10014 18760
rect 10137 18751 10195 18757
rect 10137 18717 10149 18751
rect 10183 18748 10195 18751
rect 10226 18748 10232 18760
rect 10183 18720 10232 18748
rect 10183 18717 10195 18720
rect 10137 18711 10195 18717
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 11514 18748 11520 18760
rect 10459 18720 11520 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 11514 18708 11520 18720
rect 11572 18708 11578 18760
rect 13909 18751 13967 18757
rect 12115 18717 12173 18723
rect 7193 18683 7251 18689
rect 7193 18649 7205 18683
rect 7239 18680 7251 18683
rect 8294 18680 8300 18692
rect 7239 18652 8300 18680
rect 7239 18649 7251 18652
rect 7193 18643 7251 18649
rect 8294 18640 8300 18652
rect 8352 18640 8358 18692
rect 8662 18640 8668 18692
rect 8720 18680 8726 18692
rect 9214 18680 9220 18692
rect 8720 18652 9220 18680
rect 8720 18640 8726 18652
rect 9214 18640 9220 18652
rect 9272 18640 9278 18692
rect 10772 18683 10830 18689
rect 10772 18649 10784 18683
rect 10818 18680 10830 18683
rect 11238 18680 11244 18692
rect 10818 18652 11244 18680
rect 10818 18649 10830 18652
rect 10772 18643 10830 18649
rect 11238 18640 11244 18652
rect 11296 18640 11302 18692
rect 12115 18683 12127 18717
rect 12161 18714 12173 18717
rect 13909 18717 13921 18751
rect 13955 18748 13967 18751
rect 14090 18748 14096 18760
rect 13955 18720 14096 18748
rect 13955 18717 13967 18720
rect 12161 18683 12195 18714
rect 13909 18711 13967 18717
rect 14090 18708 14096 18720
rect 14148 18708 14154 18760
rect 15396 18757 15424 18856
rect 16574 18844 16580 18856
rect 16632 18844 16638 18896
rect 17957 18887 18015 18893
rect 17957 18884 17969 18887
rect 17696 18856 17969 18884
rect 15473 18819 15531 18825
rect 15473 18785 15485 18819
rect 15519 18816 15531 18819
rect 15562 18816 15568 18828
rect 15519 18788 15568 18816
rect 15519 18785 15531 18788
rect 15473 18779 15531 18785
rect 15562 18776 15568 18788
rect 15620 18776 15626 18828
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18717 15439 18751
rect 15580 18748 15608 18776
rect 17696 18757 17724 18856
rect 17957 18853 17969 18856
rect 18003 18853 18015 18887
rect 17957 18847 18015 18853
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18104 18788 18276 18816
rect 18104 18776 18110 18788
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 15580 18720 15853 18748
rect 15381 18711 15439 18717
rect 15841 18717 15853 18720
rect 15887 18717 15899 18751
rect 15841 18711 15899 18717
rect 16669 18751 16727 18757
rect 16669 18717 16681 18751
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 17405 18751 17463 18757
rect 17405 18748 17417 18751
rect 16899 18720 17417 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 17405 18717 17417 18720
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 17681 18751 17739 18757
rect 17681 18717 17693 18751
rect 17727 18717 17739 18751
rect 17681 18711 17739 18717
rect 12115 18680 12195 18683
rect 12084 18652 12195 18680
rect 12345 18683 12403 18689
rect 12084 18624 12112 18652
rect 12345 18649 12357 18683
rect 12391 18680 12403 18683
rect 12434 18680 12440 18692
rect 12391 18652 12440 18680
rect 12391 18649 12403 18652
rect 12345 18643 12403 18649
rect 12434 18640 12440 18652
rect 12492 18680 12498 18692
rect 12618 18680 12624 18692
rect 12492 18652 12624 18680
rect 12492 18640 12498 18652
rect 12618 18640 12624 18652
rect 12676 18640 12682 18692
rect 13664 18683 13722 18689
rect 13664 18649 13676 18683
rect 13710 18680 13722 18683
rect 14366 18680 14372 18692
rect 13710 18652 14372 18680
rect 13710 18649 13722 18652
rect 13664 18643 13722 18649
rect 14366 18640 14372 18652
rect 14424 18640 14430 18692
rect 14550 18640 14556 18692
rect 14608 18680 14614 18692
rect 15194 18680 15200 18692
rect 14608 18652 15200 18680
rect 14608 18640 14614 18652
rect 15194 18640 15200 18652
rect 15252 18640 15258 18692
rect 8202 18612 8208 18624
rect 7024 18584 8208 18612
rect 8202 18572 8208 18584
rect 8260 18612 8266 18624
rect 8757 18615 8815 18621
rect 8757 18612 8769 18615
rect 8260 18584 8769 18612
rect 8260 18572 8266 18584
rect 8757 18581 8769 18584
rect 8803 18581 8815 18615
rect 8757 18575 8815 18581
rect 9953 18615 10011 18621
rect 9953 18581 9965 18615
rect 9999 18612 10011 18615
rect 10226 18612 10232 18624
rect 9999 18584 10232 18612
rect 9999 18581 10011 18584
rect 9953 18575 10011 18581
rect 10226 18572 10232 18584
rect 10284 18572 10290 18624
rect 11146 18572 11152 18624
rect 11204 18612 11210 18624
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 11204 18584 11989 18612
rect 11204 18572 11210 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 11977 18575 12035 18581
rect 12066 18572 12072 18624
rect 12124 18572 12130 18624
rect 12529 18615 12587 18621
rect 12529 18581 12541 18615
rect 12575 18612 12587 18615
rect 12802 18612 12808 18624
rect 12575 18584 12808 18612
rect 12575 18581 12587 18584
rect 12529 18575 12587 18581
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 13538 18572 13544 18624
rect 13596 18612 13602 18624
rect 15396 18612 15424 18711
rect 16684 18680 16712 18711
rect 17126 18680 17132 18692
rect 15764 18652 17132 18680
rect 15764 18621 15792 18652
rect 17126 18640 17132 18652
rect 17184 18640 17190 18692
rect 13596 18584 15424 18612
rect 15749 18615 15807 18621
rect 13596 18572 13602 18584
rect 15749 18581 15761 18615
rect 15795 18581 15807 18615
rect 17420 18612 17448 18711
rect 18138 18708 18144 18760
rect 18196 18708 18202 18760
rect 18248 18757 18276 18788
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18717 18291 18751
rect 18233 18711 18291 18717
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 20625 18751 20683 18757
rect 20625 18748 20637 18751
rect 19392 18720 20637 18748
rect 19392 18708 19398 18720
rect 20625 18717 20637 18720
rect 20671 18717 20683 18751
rect 20625 18711 20683 18717
rect 17494 18640 17500 18692
rect 17552 18680 17558 18692
rect 17957 18683 18015 18689
rect 17957 18680 17969 18683
rect 17552 18652 17969 18680
rect 17552 18640 17558 18652
rect 17957 18649 17969 18652
rect 18003 18649 18015 18683
rect 17957 18643 18015 18649
rect 18156 18612 18184 18708
rect 19886 18640 19892 18692
rect 19944 18680 19950 18692
rect 20358 18683 20416 18689
rect 20358 18680 20370 18683
rect 19944 18652 20370 18680
rect 19944 18640 19950 18652
rect 20358 18649 20370 18652
rect 20404 18649 20416 18683
rect 20358 18643 20416 18649
rect 17420 18584 18184 18612
rect 15749 18575 15807 18581
rect 19242 18572 19248 18624
rect 19300 18572 19306 18624
rect 1104 18522 22264 18544
rect 1104 18470 4255 18522
rect 4307 18470 4319 18522
rect 4371 18470 4383 18522
rect 4435 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 9545 18522
rect 9597 18470 9609 18522
rect 9661 18470 9673 18522
rect 9725 18470 9737 18522
rect 9789 18470 9801 18522
rect 9853 18470 14835 18522
rect 14887 18470 14899 18522
rect 14951 18470 14963 18522
rect 15015 18470 15027 18522
rect 15079 18470 15091 18522
rect 15143 18470 20125 18522
rect 20177 18470 20189 18522
rect 20241 18470 20253 18522
rect 20305 18470 20317 18522
rect 20369 18470 20381 18522
rect 20433 18470 22264 18522
rect 1104 18448 22264 18470
rect 2774 18368 2780 18420
rect 2832 18368 2838 18420
rect 4154 18368 4160 18420
rect 4212 18368 4218 18420
rect 4706 18408 4712 18420
rect 4448 18380 4712 18408
rect 2958 18232 2964 18284
rect 3016 18232 3022 18284
rect 4448 18281 4476 18380
rect 4706 18368 4712 18380
rect 4764 18368 4770 18420
rect 4798 18368 4804 18420
rect 4856 18368 4862 18420
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 5997 18411 6055 18417
rect 5997 18408 6009 18411
rect 5960 18380 6009 18408
rect 5960 18368 5966 18380
rect 5997 18377 6009 18380
rect 6043 18377 6055 18411
rect 5997 18371 6055 18377
rect 6362 18368 6368 18420
rect 6420 18368 6426 18420
rect 7193 18411 7251 18417
rect 7193 18377 7205 18411
rect 7239 18408 7251 18411
rect 7282 18408 7288 18420
rect 7239 18380 7288 18408
rect 7239 18377 7251 18380
rect 7193 18371 7251 18377
rect 7282 18368 7288 18380
rect 7340 18368 7346 18420
rect 8846 18368 8852 18420
rect 8904 18368 8910 18420
rect 11238 18368 11244 18420
rect 11296 18368 11302 18420
rect 11514 18368 11520 18420
rect 11572 18368 11578 18420
rect 11974 18368 11980 18420
rect 12032 18368 12038 18420
rect 13170 18368 13176 18420
rect 13228 18408 13234 18420
rect 13265 18411 13323 18417
rect 13265 18408 13277 18411
rect 13228 18380 13277 18408
rect 13228 18368 13234 18380
rect 13265 18377 13277 18380
rect 13311 18377 13323 18411
rect 13265 18371 13323 18377
rect 14366 18368 14372 18420
rect 14424 18368 14430 18420
rect 15013 18411 15071 18417
rect 15013 18377 15025 18411
rect 15059 18408 15071 18411
rect 15059 18380 15139 18408
rect 15059 18377 15071 18380
rect 15013 18371 15071 18377
rect 5074 18300 5080 18352
rect 5132 18340 5138 18352
rect 11698 18340 11704 18352
rect 5132 18312 11704 18340
rect 5132 18300 5138 18312
rect 11698 18300 11704 18312
rect 11756 18300 11762 18352
rect 4317 18275 4375 18281
rect 4317 18241 4329 18275
rect 4363 18241 4375 18275
rect 4317 18235 4375 18241
rect 4433 18275 4491 18281
rect 4433 18241 4445 18275
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 3237 18207 3295 18213
rect 3237 18173 3249 18207
rect 3283 18204 3295 18207
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 3283 18176 3433 18204
rect 3283 18173 3295 18176
rect 3237 18167 3295 18173
rect 3421 18173 3433 18176
rect 3467 18173 3479 18207
rect 3421 18167 3479 18173
rect 3970 18164 3976 18216
rect 4028 18204 4034 18216
rect 4065 18207 4123 18213
rect 4065 18204 4077 18207
rect 4028 18176 4077 18204
rect 4028 18164 4034 18176
rect 4065 18173 4077 18176
rect 4111 18204 4123 18207
rect 4347 18204 4375 18235
rect 4522 18232 4528 18284
rect 4580 18232 4586 18284
rect 4706 18232 4712 18284
rect 4764 18232 4770 18284
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18272 5043 18275
rect 5031 18244 5304 18272
rect 5031 18241 5043 18244
rect 4985 18235 5043 18241
rect 5169 18207 5227 18213
rect 5169 18204 5181 18207
rect 4111 18176 5181 18204
rect 4111 18173 4123 18176
rect 4065 18167 4123 18173
rect 5169 18173 5181 18176
rect 5215 18173 5227 18207
rect 5169 18167 5227 18173
rect 3145 18071 3203 18077
rect 3145 18037 3157 18071
rect 3191 18068 3203 18071
rect 3326 18068 3332 18080
rect 3191 18040 3332 18068
rect 3191 18037 3203 18040
rect 3145 18031 3203 18037
rect 3326 18028 3332 18040
rect 3384 18068 3390 18080
rect 5276 18068 5304 18244
rect 5534 18232 5540 18284
rect 5592 18232 5598 18284
rect 5902 18232 5908 18284
rect 5960 18232 5966 18284
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18272 6055 18275
rect 6086 18272 6092 18284
rect 6043 18244 6092 18272
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 6086 18232 6092 18244
rect 6144 18232 6150 18284
rect 6181 18275 6239 18281
rect 6181 18241 6193 18275
rect 6227 18272 6239 18275
rect 6454 18272 6460 18284
rect 6227 18244 6460 18272
rect 6227 18241 6239 18244
rect 6181 18235 6239 18241
rect 6454 18232 6460 18244
rect 6512 18232 6518 18284
rect 6546 18232 6552 18284
rect 6604 18232 6610 18284
rect 6638 18232 6644 18284
rect 6696 18272 6702 18284
rect 6917 18275 6975 18281
rect 6917 18272 6929 18275
rect 6696 18244 6929 18272
rect 6696 18232 6702 18244
rect 6917 18241 6929 18244
rect 6963 18241 6975 18275
rect 6917 18235 6975 18241
rect 7466 18232 7472 18284
rect 7524 18232 7530 18284
rect 7745 18275 7803 18281
rect 7745 18241 7757 18275
rect 7791 18241 7803 18275
rect 7745 18235 7803 18241
rect 5626 18164 5632 18216
rect 5684 18164 5690 18216
rect 5920 18204 5948 18232
rect 6733 18207 6791 18213
rect 6733 18204 6745 18207
rect 5920 18176 6745 18204
rect 6733 18173 6745 18176
rect 6779 18173 6791 18207
rect 6733 18167 6791 18173
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18173 6883 18207
rect 7484 18204 7512 18232
rect 7653 18207 7711 18213
rect 7653 18204 7665 18207
rect 7484 18176 7665 18204
rect 6825 18167 6883 18173
rect 7653 18173 7665 18176
rect 7699 18173 7711 18207
rect 7653 18167 7711 18173
rect 5905 18139 5963 18145
rect 5905 18105 5917 18139
rect 5951 18136 5963 18139
rect 5994 18136 6000 18148
rect 5951 18108 6000 18136
rect 5951 18105 5963 18108
rect 5905 18099 5963 18105
rect 5994 18096 6000 18108
rect 6052 18136 6058 18148
rect 6840 18136 6868 18167
rect 6052 18108 6868 18136
rect 6052 18096 6058 18108
rect 3384 18040 5304 18068
rect 3384 18028 3390 18040
rect 6730 18028 6736 18080
rect 6788 18068 6794 18080
rect 7760 18068 7788 18235
rect 8202 18232 8208 18284
rect 8260 18272 8266 18284
rect 8297 18275 8355 18281
rect 8297 18272 8309 18275
rect 8260 18244 8309 18272
rect 8260 18232 8266 18244
rect 8297 18241 8309 18244
rect 8343 18272 8355 18275
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 8343 18244 9229 18272
rect 8343 18241 8355 18244
rect 8297 18235 8355 18241
rect 9217 18241 9229 18244
rect 9263 18241 9275 18275
rect 9217 18235 9275 18241
rect 9944 18275 10002 18281
rect 9944 18241 9956 18275
rect 9990 18272 10002 18275
rect 10226 18272 10232 18284
rect 9990 18244 10232 18272
rect 9990 18241 10002 18244
rect 9944 18235 10002 18241
rect 10226 18232 10232 18244
rect 10284 18232 10290 18284
rect 10870 18232 10876 18284
rect 10928 18272 10934 18284
rect 11149 18275 11207 18281
rect 11149 18272 11161 18275
rect 10928 18244 11161 18272
rect 10928 18232 10934 18244
rect 11149 18241 11161 18244
rect 11195 18241 11207 18275
rect 11149 18235 11207 18241
rect 11330 18232 11336 18284
rect 11388 18232 11394 18284
rect 11992 18272 12020 18368
rect 12345 18343 12403 18349
rect 12345 18309 12357 18343
rect 12391 18340 12403 18343
rect 12618 18340 12624 18352
rect 12391 18312 12624 18340
rect 12391 18309 12403 18312
rect 12345 18303 12403 18309
rect 12618 18300 12624 18312
rect 12676 18340 12682 18352
rect 14734 18340 14740 18352
rect 12676 18312 12756 18340
rect 12676 18300 12682 18312
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 11992 18244 12265 18272
rect 12253 18241 12265 18244
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 12526 18232 12532 18284
rect 12584 18232 12590 18284
rect 12728 18281 12756 18312
rect 14292 18312 14740 18340
rect 12713 18275 12771 18281
rect 12713 18241 12725 18275
rect 12759 18241 12771 18275
rect 12713 18235 12771 18241
rect 12897 18275 12955 18281
rect 12897 18241 12909 18275
rect 12943 18272 12955 18275
rect 12986 18272 12992 18284
rect 12943 18244 12992 18272
rect 12943 18241 12955 18244
rect 12897 18235 12955 18241
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18272 13139 18275
rect 13538 18272 13544 18284
rect 13127 18244 13544 18272
rect 13127 18241 13139 18244
rect 13081 18235 13139 18241
rect 13538 18232 13544 18244
rect 13596 18232 13602 18284
rect 13722 18232 13728 18284
rect 13780 18272 13786 18284
rect 13909 18275 13967 18281
rect 13909 18272 13921 18275
rect 13780 18244 13921 18272
rect 13780 18232 13786 18244
rect 13909 18241 13921 18244
rect 13955 18241 13967 18275
rect 13909 18235 13967 18241
rect 8389 18207 8447 18213
rect 8389 18173 8401 18207
rect 8435 18173 8447 18207
rect 8389 18167 8447 18173
rect 8404 18136 8432 18167
rect 8478 18164 8484 18216
rect 8536 18204 8542 18216
rect 9125 18207 9183 18213
rect 9125 18204 9137 18207
rect 8536 18176 9137 18204
rect 8536 18164 8542 18176
rect 9125 18173 9137 18176
rect 9171 18173 9183 18207
rect 9125 18167 9183 18173
rect 9674 18164 9680 18216
rect 9732 18164 9738 18216
rect 12069 18207 12127 18213
rect 12069 18204 12081 18207
rect 11072 18176 12081 18204
rect 8570 18136 8576 18148
rect 8404 18108 8576 18136
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 9214 18096 9220 18148
rect 9272 18096 9278 18148
rect 11072 18145 11100 18176
rect 12069 18173 12081 18176
rect 12115 18204 12127 18207
rect 12434 18204 12440 18216
rect 12115 18176 12440 18204
rect 12115 18173 12127 18176
rect 12069 18167 12127 18173
rect 12434 18164 12440 18176
rect 12492 18164 12498 18216
rect 12802 18164 12808 18216
rect 12860 18204 12866 18216
rect 13740 18204 13768 18232
rect 12860 18176 13768 18204
rect 12860 18164 12866 18176
rect 13998 18164 14004 18216
rect 14056 18164 14062 18216
rect 14292 18213 14320 18312
rect 14734 18300 14740 18312
rect 14792 18300 14798 18352
rect 14918 18303 14924 18352
rect 14912 18300 14924 18303
rect 14976 18300 14982 18352
rect 14912 18297 14970 18300
rect 14553 18275 14611 18281
rect 14553 18241 14565 18275
rect 14599 18272 14611 18275
rect 14642 18272 14648 18284
rect 14599 18244 14648 18272
rect 14599 18241 14611 18244
rect 14553 18235 14611 18241
rect 14642 18232 14648 18244
rect 14700 18232 14706 18284
rect 14912 18263 14924 18297
rect 14958 18263 14970 18297
rect 14912 18257 14970 18263
rect 14277 18207 14335 18213
rect 14277 18173 14289 18207
rect 14323 18173 14335 18207
rect 14277 18167 14335 18173
rect 14826 18164 14832 18216
rect 14884 18204 14890 18216
rect 15111 18204 15139 18380
rect 15194 18300 15200 18352
rect 15252 18340 15258 18352
rect 17494 18340 17500 18352
rect 15252 18312 17500 18340
rect 15252 18300 15258 18312
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 16853 18275 16911 18281
rect 16853 18241 16865 18275
rect 16899 18241 16911 18275
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 16853 18235 16911 18241
rect 17052 18244 17233 18272
rect 14884 18176 15139 18204
rect 14884 18164 14890 18176
rect 11057 18139 11115 18145
rect 11057 18105 11069 18139
rect 11103 18105 11115 18139
rect 11057 18099 11115 18105
rect 14642 18096 14648 18148
rect 14700 18136 14706 18148
rect 15197 18139 15255 18145
rect 15197 18136 15209 18139
rect 14700 18108 15209 18136
rect 14700 18096 14706 18108
rect 15197 18105 15209 18108
rect 15243 18105 15255 18139
rect 16868 18136 16896 18235
rect 17052 18216 17080 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18241 17371 18275
rect 17313 18235 17371 18241
rect 17034 18164 17040 18216
rect 17092 18164 17098 18216
rect 17126 18164 17132 18216
rect 17184 18204 17190 18216
rect 17328 18204 17356 18235
rect 17184 18176 17356 18204
rect 17184 18164 17190 18176
rect 17497 18139 17555 18145
rect 17497 18136 17509 18139
rect 16868 18108 17509 18136
rect 15197 18099 15255 18105
rect 17497 18105 17509 18108
rect 17543 18105 17555 18139
rect 17497 18099 17555 18105
rect 6788 18040 7788 18068
rect 6788 18028 6794 18040
rect 8754 18028 8760 18080
rect 8812 18068 8818 18080
rect 9232 18068 9260 18096
rect 14550 18068 14556 18080
rect 8812 18040 14556 18068
rect 8812 18028 8818 18040
rect 14550 18028 14556 18040
rect 14608 18028 14614 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 14918 18068 14924 18080
rect 14792 18040 14924 18068
rect 14792 18028 14798 18040
rect 14918 18028 14924 18040
rect 14976 18028 14982 18080
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 16669 18071 16727 18077
rect 16669 18068 16681 18071
rect 16632 18040 16681 18068
rect 16632 18028 16638 18040
rect 16669 18037 16681 18040
rect 16715 18037 16727 18071
rect 16669 18031 16727 18037
rect 17034 18028 17040 18080
rect 17092 18028 17098 18080
rect 1104 17978 22264 18000
rect 1104 17926 3595 17978
rect 3647 17926 3659 17978
rect 3711 17926 3723 17978
rect 3775 17926 3787 17978
rect 3839 17926 3851 17978
rect 3903 17926 8885 17978
rect 8937 17926 8949 17978
rect 9001 17926 9013 17978
rect 9065 17926 9077 17978
rect 9129 17926 9141 17978
rect 9193 17926 14175 17978
rect 14227 17926 14239 17978
rect 14291 17926 14303 17978
rect 14355 17926 14367 17978
rect 14419 17926 14431 17978
rect 14483 17926 19465 17978
rect 19517 17926 19529 17978
rect 19581 17926 19593 17978
rect 19645 17926 19657 17978
rect 19709 17926 19721 17978
rect 19773 17926 22264 17978
rect 1104 17904 22264 17926
rect 9950 17824 9956 17876
rect 10008 17864 10014 17876
rect 10413 17867 10471 17873
rect 10413 17864 10425 17867
rect 10008 17836 10425 17864
rect 10008 17824 10014 17836
rect 10413 17833 10425 17836
rect 10459 17833 10471 17867
rect 10413 17827 10471 17833
rect 11330 17824 11336 17876
rect 11388 17864 11394 17876
rect 12069 17867 12127 17873
rect 12069 17864 12081 17867
rect 11388 17836 12081 17864
rect 11388 17824 11394 17836
rect 12069 17833 12081 17836
rect 12115 17833 12127 17867
rect 12069 17827 12127 17833
rect 12250 17824 12256 17876
rect 12308 17824 12314 17876
rect 14461 17867 14519 17873
rect 14461 17833 14473 17867
rect 14507 17864 14519 17867
rect 16022 17864 16028 17876
rect 14507 17836 16028 17864
rect 14507 17833 14519 17836
rect 14461 17827 14519 17833
rect 16022 17824 16028 17836
rect 16080 17824 16086 17876
rect 16117 17867 16175 17873
rect 16117 17833 16129 17867
rect 16163 17864 16175 17867
rect 17034 17864 17040 17876
rect 16163 17836 17040 17864
rect 16163 17833 16175 17836
rect 16117 17827 16175 17833
rect 17034 17824 17040 17836
rect 17092 17824 17098 17876
rect 17402 17824 17408 17876
rect 17460 17864 17466 17876
rect 17681 17867 17739 17873
rect 17681 17864 17693 17867
rect 17460 17836 17693 17864
rect 17460 17824 17466 17836
rect 17681 17833 17693 17836
rect 17727 17833 17739 17867
rect 17681 17827 17739 17833
rect 10321 17799 10379 17805
rect 10321 17765 10333 17799
rect 10367 17796 10379 17799
rect 10367 17768 11008 17796
rect 10367 17765 10379 17768
rect 10321 17759 10379 17765
rect 4062 17688 4068 17740
rect 4120 17728 4126 17740
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 4120 17700 4445 17728
rect 4120 17688 4126 17700
rect 4433 17697 4445 17700
rect 4479 17728 4491 17731
rect 4522 17728 4528 17740
rect 4479 17700 4528 17728
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 4522 17688 4528 17700
rect 4580 17688 4586 17740
rect 10980 17737 11008 17768
rect 10965 17731 11023 17737
rect 9968 17700 10180 17728
rect 3326 17620 3332 17672
rect 3384 17660 3390 17672
rect 3421 17663 3479 17669
rect 3421 17660 3433 17663
rect 3384 17632 3433 17660
rect 3384 17620 3390 17632
rect 3421 17629 3433 17632
rect 3467 17629 3479 17663
rect 3421 17623 3479 17629
rect 3510 17620 3516 17672
rect 3568 17660 3574 17672
rect 3605 17663 3663 17669
rect 3605 17660 3617 17663
rect 3568 17632 3617 17660
rect 3568 17620 3574 17632
rect 3605 17629 3617 17632
rect 3651 17629 3663 17663
rect 3605 17623 3663 17629
rect 4985 17663 5043 17669
rect 4985 17629 4997 17663
rect 5031 17660 5043 17663
rect 5534 17660 5540 17672
rect 5031 17632 5540 17660
rect 5031 17629 5043 17632
rect 4985 17623 5043 17629
rect 3620 17592 3648 17623
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 9306 17620 9312 17672
rect 9364 17660 9370 17672
rect 9968 17669 9996 17700
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9364 17632 9781 17660
rect 9364 17620 9370 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9769 17623 9827 17629
rect 9953 17663 10011 17669
rect 9953 17629 9965 17663
rect 9999 17629 10011 17663
rect 9953 17623 10011 17629
rect 10042 17620 10048 17672
rect 10100 17620 10106 17672
rect 10152 17660 10180 17700
rect 10965 17697 10977 17731
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 12161 17731 12219 17737
rect 12161 17697 12173 17731
rect 12207 17728 12219 17731
rect 12268 17728 12296 17824
rect 13722 17756 13728 17808
rect 13780 17796 13786 17808
rect 13780 17768 15608 17796
rect 13780 17756 13786 17768
rect 13740 17728 13768 17756
rect 14826 17728 14832 17740
rect 12207 17700 12296 17728
rect 12728 17700 13768 17728
rect 14661 17700 14832 17728
rect 12207 17697 12219 17700
rect 12161 17691 12219 17697
rect 10152 17632 11192 17660
rect 3620 17564 5212 17592
rect 5184 17536 5212 17564
rect 10318 17552 10324 17604
rect 10376 17552 10382 17604
rect 11164 17601 11192 17632
rect 11330 17620 11336 17672
rect 11388 17660 11394 17672
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 11388 17632 11713 17660
rect 11388 17620 11394 17632
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11701 17623 11759 17629
rect 11882 17620 11888 17672
rect 11940 17620 11946 17672
rect 11977 17663 12035 17669
rect 11977 17629 11989 17663
rect 12023 17660 12035 17663
rect 12066 17660 12072 17672
rect 12023 17632 12072 17660
rect 12023 17629 12035 17632
rect 11977 17623 12035 17629
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 12618 17620 12624 17672
rect 12676 17620 12682 17672
rect 12728 17669 12756 17700
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17629 12771 17663
rect 12713 17623 12771 17629
rect 12989 17663 13047 17669
rect 12989 17629 13001 17663
rect 13035 17660 13047 17663
rect 13446 17660 13452 17672
rect 13035 17632 13452 17660
rect 13035 17629 13047 17632
rect 12989 17623 13047 17629
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 14661 17669 14689 17700
rect 14826 17688 14832 17700
rect 14884 17688 14890 17740
rect 15580 17737 15608 17768
rect 15197 17731 15255 17737
rect 15197 17728 15209 17731
rect 15028 17700 15209 17728
rect 15028 17669 15056 17700
rect 15197 17697 15209 17700
rect 15243 17697 15255 17731
rect 15197 17691 15255 17697
rect 15565 17731 15623 17737
rect 15565 17697 15577 17731
rect 15611 17697 15623 17731
rect 15565 17691 15623 17697
rect 14645 17663 14703 17669
rect 14645 17629 14657 17663
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17629 15071 17663
rect 15013 17623 15071 17629
rect 15105 17663 15163 17669
rect 15105 17629 15117 17663
rect 15151 17660 15163 17663
rect 15286 17660 15292 17672
rect 15151 17632 15292 17660
rect 15151 17629 15163 17632
rect 15105 17623 15163 17629
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 16040 17669 16068 17824
rect 15381 17663 15439 17669
rect 15381 17629 15393 17663
rect 15427 17629 15439 17663
rect 15381 17623 15439 17629
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17629 16083 17663
rect 16025 17623 16083 17629
rect 11149 17595 11207 17601
rect 11149 17561 11161 17595
rect 11195 17592 11207 17595
rect 12805 17595 12863 17601
rect 11195 17564 12664 17592
rect 11195 17561 11207 17564
rect 11149 17555 11207 17561
rect 3510 17484 3516 17536
rect 3568 17484 3574 17536
rect 3786 17484 3792 17536
rect 3844 17484 3850 17536
rect 4154 17484 4160 17536
rect 4212 17524 4218 17536
rect 4706 17524 4712 17536
rect 4212 17496 4712 17524
rect 4212 17484 4218 17496
rect 4706 17484 4712 17496
rect 4764 17524 4770 17536
rect 4893 17527 4951 17533
rect 4893 17524 4905 17527
rect 4764 17496 4905 17524
rect 4764 17484 4770 17496
rect 4893 17493 4905 17496
rect 4939 17493 4951 17527
rect 4893 17487 4951 17493
rect 5166 17484 5172 17536
rect 5224 17484 5230 17536
rect 9306 17484 9312 17536
rect 9364 17524 9370 17536
rect 9861 17527 9919 17533
rect 9861 17524 9873 17527
rect 9364 17496 9873 17524
rect 9364 17484 9370 17496
rect 9861 17493 9873 17496
rect 9907 17493 9919 17527
rect 9861 17487 9919 17493
rect 10134 17484 10140 17536
rect 10192 17484 10198 17536
rect 12434 17484 12440 17536
rect 12492 17484 12498 17536
rect 12636 17524 12664 17564
rect 12805 17561 12817 17595
rect 12851 17592 12863 17595
rect 13262 17592 13268 17604
rect 12851 17564 13268 17592
rect 12851 17561 12863 17564
rect 12805 17555 12863 17561
rect 13262 17552 13268 17564
rect 13320 17552 13326 17604
rect 14550 17552 14556 17604
rect 14608 17592 14614 17604
rect 14737 17595 14795 17601
rect 14737 17592 14749 17595
rect 14608 17564 14749 17592
rect 14608 17552 14614 17564
rect 14737 17561 14749 17564
rect 14783 17561 14795 17595
rect 14737 17555 14795 17561
rect 14829 17595 14887 17601
rect 14829 17561 14841 17595
rect 14875 17561 14887 17595
rect 15396 17592 15424 17623
rect 16206 17620 16212 17672
rect 16264 17620 16270 17672
rect 16574 17669 16580 17672
rect 16301 17663 16359 17669
rect 16301 17629 16313 17663
rect 16347 17629 16359 17663
rect 16568 17660 16580 17669
rect 16535 17632 16580 17660
rect 16301 17623 16359 17629
rect 16568 17623 16580 17632
rect 16316 17592 16344 17623
rect 16574 17620 16580 17623
rect 16632 17620 16638 17672
rect 16942 17620 16948 17672
rect 17000 17620 17006 17672
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 19794 17660 19800 17672
rect 19751 17632 19800 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 19794 17620 19800 17632
rect 19852 17620 19858 17672
rect 21450 17620 21456 17672
rect 21508 17620 21514 17672
rect 16960 17592 16988 17620
rect 15396 17564 15608 17592
rect 16316 17564 16988 17592
rect 14829 17555 14887 17561
rect 12986 17524 12992 17536
rect 12636 17496 12992 17524
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 14642 17484 14648 17536
rect 14700 17524 14706 17536
rect 14844 17524 14872 17555
rect 15580 17536 15608 17564
rect 14700 17496 14872 17524
rect 14700 17484 14706 17496
rect 15562 17484 15568 17536
rect 15620 17484 15626 17536
rect 19886 17484 19892 17536
rect 19944 17484 19950 17536
rect 20898 17484 20904 17536
rect 20956 17484 20962 17536
rect 1104 17434 22264 17456
rect 1104 17382 4255 17434
rect 4307 17382 4319 17434
rect 4371 17382 4383 17434
rect 4435 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 9545 17434
rect 9597 17382 9609 17434
rect 9661 17382 9673 17434
rect 9725 17382 9737 17434
rect 9789 17382 9801 17434
rect 9853 17382 14835 17434
rect 14887 17382 14899 17434
rect 14951 17382 14963 17434
rect 15015 17382 15027 17434
rect 15079 17382 15091 17434
rect 15143 17382 20125 17434
rect 20177 17382 20189 17434
rect 20241 17382 20253 17434
rect 20305 17382 20317 17434
rect 20369 17382 20381 17434
rect 20433 17382 22264 17434
rect 1104 17360 22264 17382
rect 3510 17280 3516 17332
rect 3568 17280 3574 17332
rect 3786 17280 3792 17332
rect 3844 17280 3850 17332
rect 3881 17323 3939 17329
rect 3881 17289 3893 17323
rect 3927 17320 3939 17323
rect 4614 17320 4620 17332
rect 3927 17292 4620 17320
rect 3927 17289 3939 17292
rect 3881 17283 3939 17289
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 10318 17280 10324 17332
rect 10376 17320 10382 17332
rect 10689 17323 10747 17329
rect 10689 17320 10701 17323
rect 10376 17292 10701 17320
rect 10376 17280 10382 17292
rect 10689 17289 10701 17292
rect 10735 17289 10747 17323
rect 10689 17283 10747 17289
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12526 17320 12532 17332
rect 12483 17292 12532 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 14642 17280 14648 17332
rect 14700 17280 14706 17332
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 15105 17323 15163 17329
rect 15105 17320 15117 17323
rect 14792 17292 15117 17320
rect 14792 17280 14798 17292
rect 15105 17289 15117 17292
rect 15151 17289 15163 17323
rect 15105 17283 15163 17289
rect 19886 17280 19892 17332
rect 19944 17280 19950 17332
rect 21269 17323 21327 17329
rect 21269 17289 21281 17323
rect 21315 17320 21327 17323
rect 21450 17320 21456 17332
rect 21315 17292 21456 17320
rect 21315 17289 21327 17292
rect 21269 17283 21327 17289
rect 21450 17280 21456 17292
rect 21508 17280 21514 17332
rect 1397 17187 1455 17193
rect 1397 17153 1409 17187
rect 1443 17184 1455 17187
rect 1486 17184 1492 17196
rect 1443 17156 1492 17184
rect 1443 17153 1455 17156
rect 1397 17147 1455 17153
rect 1486 17144 1492 17156
rect 1544 17144 1550 17196
rect 1664 17187 1722 17193
rect 1664 17153 1676 17187
rect 1710 17184 1722 17187
rect 2869 17187 2927 17193
rect 2869 17184 2881 17187
rect 1710 17156 2881 17184
rect 1710 17153 1722 17156
rect 1664 17147 1722 17153
rect 2869 17153 2881 17156
rect 2915 17153 2927 17187
rect 2869 17147 2927 17153
rect 3053 17187 3111 17193
rect 3053 17153 3065 17187
rect 3099 17184 3111 17187
rect 3528 17184 3556 17280
rect 3099 17156 3556 17184
rect 3099 17153 3111 17156
rect 3053 17147 3111 17153
rect 3602 17144 3608 17196
rect 3660 17144 3666 17196
rect 3804 17184 3832 17280
rect 3712 17156 3832 17184
rect 3988 17224 4476 17252
rect 3329 17119 3387 17125
rect 3329 17085 3341 17119
rect 3375 17116 3387 17119
rect 3712 17116 3740 17156
rect 3375 17088 3740 17116
rect 3789 17119 3847 17125
rect 3375 17085 3387 17088
rect 3329 17079 3387 17085
rect 3789 17085 3801 17119
rect 3835 17116 3847 17119
rect 3988 17116 4016 17224
rect 4448 17196 4476 17224
rect 6178 17212 6184 17264
rect 6236 17252 6242 17264
rect 6365 17255 6423 17261
rect 6365 17252 6377 17255
rect 6236 17224 6377 17252
rect 6236 17212 6242 17224
rect 6365 17221 6377 17224
rect 6411 17221 6423 17255
rect 6365 17215 6423 17221
rect 9490 17212 9496 17264
rect 9548 17252 9554 17264
rect 13906 17252 13912 17264
rect 9548 17224 13912 17252
rect 9548 17212 9554 17224
rect 13906 17212 13912 17224
rect 13964 17212 13970 17264
rect 14550 17212 14556 17264
rect 14608 17212 14614 17264
rect 14660 17252 14688 17280
rect 15197 17255 15255 17261
rect 15197 17252 15209 17255
rect 14660 17224 15209 17252
rect 4065 17187 4123 17193
rect 4065 17153 4077 17187
rect 4111 17184 4123 17187
rect 4154 17184 4160 17196
rect 4111 17156 4160 17184
rect 4111 17153 4123 17156
rect 4065 17147 4123 17153
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4430 17144 4436 17196
rect 4488 17144 4494 17196
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17184 4675 17187
rect 4706 17184 4712 17196
rect 4663 17156 4712 17184
rect 4663 17153 4675 17156
rect 4617 17147 4675 17153
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 5626 17144 5632 17196
rect 5684 17144 5690 17196
rect 6546 17144 6552 17196
rect 6604 17144 6610 17196
rect 6638 17144 6644 17196
rect 6696 17144 6702 17196
rect 7282 17144 7288 17196
rect 7340 17144 7346 17196
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17184 7527 17187
rect 7834 17184 7840 17196
rect 7515 17156 7840 17184
rect 7515 17153 7527 17156
rect 7469 17147 7527 17153
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 9306 17193 9312 17196
rect 8297 17187 8355 17193
rect 8297 17153 8309 17187
rect 8343 17153 8355 17187
rect 8297 17147 8355 17153
rect 9289 17187 9312 17193
rect 9289 17153 9301 17187
rect 9289 17147 9312 17153
rect 3835 17088 4016 17116
rect 4249 17119 4307 17125
rect 3835 17085 3847 17088
rect 3789 17079 3847 17085
rect 4249 17085 4261 17119
rect 4295 17085 4307 17119
rect 4249 17079 4307 17085
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17116 4399 17119
rect 4387 17088 5304 17116
rect 4387 17085 4399 17088
rect 4341 17079 4399 17085
rect 2777 17051 2835 17057
rect 2777 17017 2789 17051
rect 2823 17048 2835 17051
rect 4062 17048 4068 17060
rect 2823 17020 4068 17048
rect 2823 17017 2835 17020
rect 2777 17011 2835 17017
rect 4062 17008 4068 17020
rect 4120 17048 4126 17060
rect 4264 17048 4292 17079
rect 4120 17020 4292 17048
rect 4120 17008 4126 17020
rect 5276 16992 5304 17088
rect 7098 17076 7104 17128
rect 7156 17116 7162 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7156 17088 8033 17116
rect 7156 17076 7162 17088
rect 8021 17085 8033 17088
rect 8067 17116 8079 17119
rect 8113 17119 8171 17125
rect 8113 17116 8125 17119
rect 8067 17088 8125 17116
rect 8067 17085 8079 17088
rect 8021 17079 8079 17085
rect 8113 17085 8125 17088
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 7745 17051 7803 17057
rect 7745 17017 7757 17051
rect 7791 17048 7803 17051
rect 8202 17048 8208 17060
rect 7791 17020 8208 17048
rect 7791 17017 7803 17020
rect 7745 17011 7803 17017
rect 8202 17008 8208 17020
rect 8260 17008 8266 17060
rect 8312 17048 8340 17147
rect 9306 17144 9312 17147
rect 9364 17144 9370 17196
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 8481 17119 8539 17125
rect 8481 17085 8493 17119
rect 8527 17116 8539 17119
rect 8570 17116 8576 17128
rect 8527 17088 8576 17116
rect 8527 17085 8539 17088
rect 8481 17079 8539 17085
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 9033 17119 9091 17125
rect 9033 17085 9045 17119
rect 9079 17085 9091 17119
rect 9033 17079 9091 17085
rect 8312 17020 8524 17048
rect 8496 16992 8524 17020
rect 3234 16940 3240 16992
rect 3292 16980 3298 16992
rect 3421 16983 3479 16989
rect 3421 16980 3433 16983
rect 3292 16952 3433 16980
rect 3292 16940 3298 16952
rect 3421 16949 3433 16952
rect 3467 16949 3479 16983
rect 3421 16943 3479 16949
rect 5258 16940 5264 16992
rect 5316 16980 5322 16992
rect 5537 16983 5595 16989
rect 5537 16980 5549 16983
rect 5316 16952 5549 16980
rect 5316 16940 5322 16952
rect 5537 16949 5549 16952
rect 5583 16949 5595 16983
rect 5537 16943 5595 16949
rect 6086 16940 6092 16992
rect 6144 16980 6150 16992
rect 6365 16983 6423 16989
rect 6365 16980 6377 16983
rect 6144 16952 6377 16980
rect 6144 16940 6150 16952
rect 6365 16949 6377 16952
rect 6411 16949 6423 16983
rect 6365 16943 6423 16949
rect 7466 16940 7472 16992
rect 7524 16940 7530 16992
rect 7558 16940 7564 16992
rect 7616 16940 7622 16992
rect 8478 16940 8484 16992
rect 8536 16940 8542 16992
rect 9048 16980 9076 17079
rect 11238 17076 11244 17128
rect 11296 17076 11302 17128
rect 11609 17119 11667 17125
rect 11609 17085 11621 17119
rect 11655 17116 11667 17119
rect 12250 17116 12256 17128
rect 11655 17088 12256 17116
rect 11655 17085 11667 17088
rect 11609 17079 11667 17085
rect 12250 17076 12256 17088
rect 12308 17076 12314 17128
rect 12526 17076 12532 17128
rect 12584 17116 12590 17128
rect 12636 17116 12664 17147
rect 12802 17144 12808 17196
rect 12860 17144 12866 17196
rect 12894 17144 12900 17196
rect 12952 17144 12958 17196
rect 12986 17144 12992 17196
rect 13044 17144 13050 17196
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17153 13323 17187
rect 13265 17147 13323 17153
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17153 14519 17187
rect 14461 17147 14519 17153
rect 12584 17088 12664 17116
rect 12584 17076 12590 17088
rect 13280 17048 13308 17147
rect 12406 17020 13308 17048
rect 14476 17048 14504 17147
rect 14568 17116 14596 17212
rect 14660 17193 14688 17224
rect 15197 17221 15209 17224
rect 15243 17221 15255 17255
rect 15197 17215 15255 17221
rect 15562 17212 15568 17264
rect 15620 17212 15626 17264
rect 19334 17252 19340 17264
rect 18432 17224 19340 17252
rect 14645 17187 14703 17193
rect 14645 17153 14657 17187
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 14737 17187 14795 17193
rect 14737 17153 14749 17187
rect 14783 17153 14795 17187
rect 14737 17147 14795 17153
rect 14829 17187 14887 17193
rect 14829 17153 14841 17187
rect 14875 17184 14887 17187
rect 15286 17184 15292 17196
rect 14875 17156 15292 17184
rect 14875 17153 14887 17156
rect 14829 17147 14887 17153
rect 14752 17116 14780 17147
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17184 15439 17187
rect 15470 17184 15476 17196
rect 15427 17156 15476 17184
rect 15427 17153 15439 17156
rect 15381 17147 15439 17153
rect 15470 17144 15476 17156
rect 15528 17144 15534 17196
rect 16206 17144 16212 17196
rect 16264 17144 16270 17196
rect 14568 17088 14780 17116
rect 15194 17048 15200 17060
rect 14476 17020 15200 17048
rect 9398 16980 9404 16992
rect 9048 16952 9404 16980
rect 9398 16940 9404 16952
rect 9456 16940 9462 16992
rect 10042 16940 10048 16992
rect 10100 16980 10106 16992
rect 10413 16983 10471 16989
rect 10413 16980 10425 16983
rect 10100 16952 10425 16980
rect 10100 16940 10106 16952
rect 10413 16949 10425 16952
rect 10459 16980 10471 16983
rect 11330 16980 11336 16992
rect 10459 16952 11336 16980
rect 10459 16949 10471 16952
rect 10413 16943 10471 16949
rect 11330 16940 11336 16952
rect 11388 16940 11394 16992
rect 11606 16940 11612 16992
rect 11664 16980 11670 16992
rect 12161 16983 12219 16989
rect 12161 16980 12173 16983
rect 11664 16952 12173 16980
rect 11664 16940 11670 16952
rect 12161 16949 12173 16952
rect 12207 16980 12219 16983
rect 12406 16980 12434 17020
rect 15194 17008 15200 17020
rect 15252 17048 15258 17060
rect 16224 17048 16252 17144
rect 16942 17076 16948 17128
rect 17000 17116 17006 17128
rect 18432 17125 18460 17224
rect 19334 17212 19340 17224
rect 19392 17212 19398 17264
rect 19904 17252 19932 17280
rect 20134 17255 20192 17261
rect 20134 17252 20146 17255
rect 19904 17224 20146 17252
rect 20134 17221 20146 17224
rect 20180 17221 20192 17255
rect 20134 17215 20192 17221
rect 18506 17144 18512 17196
rect 18564 17184 18570 17196
rect 18673 17187 18731 17193
rect 18673 17184 18685 17187
rect 18564 17156 18685 17184
rect 18564 17144 18570 17156
rect 18673 17153 18685 17156
rect 18719 17153 18731 17187
rect 19352 17184 19380 17212
rect 19886 17184 19892 17196
rect 19352 17156 19892 17184
rect 18673 17147 18731 17153
rect 19886 17144 19892 17156
rect 19944 17144 19950 17196
rect 18417 17119 18475 17125
rect 18417 17116 18429 17119
rect 17000 17088 18429 17116
rect 17000 17076 17006 17088
rect 18417 17085 18429 17088
rect 18463 17085 18475 17119
rect 18417 17079 18475 17085
rect 15252 17020 16252 17048
rect 15252 17008 15258 17020
rect 12207 16952 12434 16980
rect 12207 16949 12219 16952
rect 12161 16943 12219 16949
rect 12986 16940 12992 16992
rect 13044 16980 13050 16992
rect 13081 16983 13139 16989
rect 13081 16980 13093 16983
rect 13044 16952 13093 16980
rect 13044 16940 13050 16952
rect 13081 16949 13093 16952
rect 13127 16949 13139 16983
rect 13081 16943 13139 16949
rect 13354 16940 13360 16992
rect 13412 16940 13418 16992
rect 19797 16983 19855 16989
rect 19797 16949 19809 16983
rect 19843 16980 19855 16983
rect 20070 16980 20076 16992
rect 19843 16952 20076 16980
rect 19843 16949 19855 16952
rect 19797 16943 19855 16949
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 1104 16890 22264 16912
rect 1104 16838 3595 16890
rect 3647 16838 3659 16890
rect 3711 16838 3723 16890
rect 3775 16838 3787 16890
rect 3839 16838 3851 16890
rect 3903 16838 8885 16890
rect 8937 16838 8949 16890
rect 9001 16838 9013 16890
rect 9065 16838 9077 16890
rect 9129 16838 9141 16890
rect 9193 16838 14175 16890
rect 14227 16838 14239 16890
rect 14291 16838 14303 16890
rect 14355 16838 14367 16890
rect 14419 16838 14431 16890
rect 14483 16838 19465 16890
rect 19517 16838 19529 16890
rect 19581 16838 19593 16890
rect 19645 16838 19657 16890
rect 19709 16838 19721 16890
rect 19773 16838 22264 16890
rect 1104 16816 22264 16838
rect 3053 16779 3111 16785
rect 3053 16745 3065 16779
rect 3099 16776 3111 16779
rect 3421 16779 3479 16785
rect 3421 16776 3433 16779
rect 3099 16748 3433 16776
rect 3099 16745 3111 16748
rect 3053 16739 3111 16745
rect 3421 16745 3433 16748
rect 3467 16776 3479 16779
rect 4890 16776 4896 16788
rect 3467 16748 4476 16776
rect 3467 16745 3479 16748
rect 3421 16739 3479 16745
rect 3237 16711 3295 16717
rect 3237 16677 3249 16711
rect 3283 16708 3295 16711
rect 3326 16708 3332 16720
rect 3283 16680 3332 16708
rect 3283 16677 3295 16680
rect 3237 16671 3295 16677
rect 3326 16668 3332 16680
rect 3384 16668 3390 16720
rect 1486 16600 1492 16652
rect 1544 16640 1550 16652
rect 1673 16643 1731 16649
rect 1673 16640 1685 16643
rect 1544 16612 1685 16640
rect 1544 16600 1550 16612
rect 1673 16609 1685 16612
rect 1719 16640 1731 16643
rect 1719 16612 1753 16640
rect 1719 16609 1731 16612
rect 1673 16603 1731 16609
rect 1688 16448 1716 16603
rect 4448 16584 4476 16748
rect 4632 16748 4896 16776
rect 4632 16652 4660 16748
rect 4890 16736 4896 16748
rect 4948 16736 4954 16788
rect 5626 16736 5632 16788
rect 5684 16776 5690 16788
rect 5997 16779 6055 16785
rect 5997 16776 6009 16779
rect 5684 16748 6009 16776
rect 5684 16736 5690 16748
rect 5997 16745 6009 16748
rect 6043 16776 6055 16779
rect 6362 16776 6368 16788
rect 6043 16748 6368 16776
rect 6043 16745 6055 16748
rect 5997 16739 6055 16745
rect 6362 16736 6368 16748
rect 6420 16736 6426 16788
rect 6454 16736 6460 16788
rect 6512 16736 6518 16788
rect 7374 16776 7380 16788
rect 7208 16748 7380 16776
rect 7098 16668 7104 16720
rect 7156 16668 7162 16720
rect 4614 16600 4620 16652
rect 4672 16600 4678 16652
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 6604 16612 6684 16640
rect 6604 16600 6610 16612
rect 3510 16532 3516 16584
rect 3568 16532 3574 16584
rect 4430 16532 4436 16584
rect 4488 16572 4494 16584
rect 6656 16581 6684 16612
rect 6641 16575 6699 16581
rect 4488 16544 4844 16572
rect 4488 16532 4494 16544
rect 1940 16507 1998 16513
rect 1940 16473 1952 16507
rect 1986 16504 1998 16507
rect 2130 16504 2136 16516
rect 1986 16476 2136 16504
rect 1986 16473 1998 16476
rect 1940 16467 1998 16473
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 3405 16507 3463 16513
rect 3405 16473 3417 16507
rect 3451 16504 3463 16507
rect 3528 16504 3556 16532
rect 3451 16476 3556 16504
rect 3605 16507 3663 16513
rect 3451 16473 3463 16476
rect 3405 16467 3463 16473
rect 3605 16473 3617 16507
rect 3651 16504 3663 16507
rect 4062 16504 4068 16516
rect 3651 16476 4068 16504
rect 3651 16473 3663 16476
rect 3605 16467 3663 16473
rect 4062 16464 4068 16476
rect 4120 16464 4126 16516
rect 4816 16448 4844 16544
rect 6641 16541 6653 16575
rect 6687 16541 6699 16575
rect 6641 16535 6699 16541
rect 6914 16532 6920 16584
rect 6972 16532 6978 16584
rect 7116 16581 7144 16668
rect 7208 16649 7236 16748
rect 7374 16736 7380 16748
rect 7432 16776 7438 16788
rect 12066 16776 12072 16788
rect 7432 16748 9444 16776
rect 7432 16736 7438 16748
rect 8202 16668 8208 16720
rect 8260 16708 8266 16720
rect 8941 16711 8999 16717
rect 8941 16708 8953 16711
rect 8260 16680 8953 16708
rect 8260 16668 8266 16680
rect 8941 16677 8953 16680
rect 8987 16677 8999 16711
rect 8941 16671 8999 16677
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16609 7251 16643
rect 7193 16603 7251 16609
rect 7466 16581 7472 16584
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16541 7159 16575
rect 7460 16572 7472 16581
rect 7427 16544 7472 16572
rect 7101 16535 7159 16541
rect 7460 16535 7472 16544
rect 7466 16532 7472 16535
rect 7524 16532 7530 16584
rect 4884 16507 4942 16513
rect 4884 16473 4896 16507
rect 4930 16504 4942 16507
rect 5718 16504 5724 16516
rect 4930 16476 5724 16504
rect 4930 16473 4942 16476
rect 4884 16467 4942 16473
rect 5718 16464 5724 16476
rect 5776 16464 5782 16516
rect 6733 16507 6791 16513
rect 6733 16473 6745 16507
rect 6779 16473 6791 16507
rect 6733 16467 6791 16473
rect 6825 16507 6883 16513
rect 6825 16473 6837 16507
rect 6871 16504 6883 16507
rect 8220 16504 8248 16668
rect 9416 16652 9444 16748
rect 9692 16748 12072 16776
rect 9692 16717 9720 16748
rect 12066 16736 12072 16748
rect 12124 16736 12130 16788
rect 12802 16736 12808 16788
rect 12860 16736 12866 16788
rect 12894 16736 12900 16788
rect 12952 16736 12958 16788
rect 14642 16736 14648 16788
rect 14700 16736 14706 16788
rect 15286 16736 15292 16788
rect 15344 16776 15350 16788
rect 15381 16779 15439 16785
rect 15381 16776 15393 16779
rect 15344 16748 15393 16776
rect 15344 16736 15350 16748
rect 15381 16745 15393 16748
rect 15427 16745 15439 16779
rect 15381 16739 15439 16745
rect 17865 16779 17923 16785
rect 17865 16745 17877 16779
rect 17911 16776 17923 16779
rect 18506 16776 18512 16788
rect 17911 16748 18512 16776
rect 17911 16745 17923 16748
rect 17865 16739 17923 16745
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 19705 16779 19763 16785
rect 19705 16745 19717 16779
rect 19751 16776 19763 16779
rect 19794 16776 19800 16788
rect 19751 16748 19800 16776
rect 19751 16745 19763 16748
rect 19705 16739 19763 16745
rect 19794 16736 19800 16748
rect 19852 16736 19858 16788
rect 20898 16736 20904 16788
rect 20956 16736 20962 16788
rect 9677 16711 9735 16717
rect 9677 16677 9689 16711
rect 9723 16677 9735 16711
rect 9677 16671 9735 16677
rect 11238 16668 11244 16720
rect 11296 16708 11302 16720
rect 12618 16708 12624 16720
rect 11296 16680 12624 16708
rect 11296 16668 11302 16680
rect 12618 16668 12624 16680
rect 12676 16668 12682 16720
rect 14660 16708 14688 16736
rect 14921 16711 14979 16717
rect 14921 16708 14933 16711
rect 14660 16680 14933 16708
rect 14921 16677 14933 16680
rect 14967 16677 14979 16711
rect 14921 16671 14979 16677
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 9456 16612 9873 16640
rect 9456 16600 9462 16612
rect 9861 16609 9873 16612
rect 9907 16609 9919 16643
rect 9861 16603 9919 16609
rect 11977 16643 12035 16649
rect 11977 16609 11989 16643
rect 12023 16640 12035 16643
rect 12434 16640 12440 16652
rect 12023 16612 12440 16640
rect 12023 16609 12035 16612
rect 11977 16603 12035 16609
rect 9309 16575 9367 16581
rect 9309 16572 9321 16575
rect 8496 16544 9321 16572
rect 8496 16516 8524 16544
rect 9309 16541 9321 16544
rect 9355 16541 9367 16575
rect 9309 16535 9367 16541
rect 9490 16532 9496 16584
rect 9548 16532 9554 16584
rect 9766 16532 9772 16584
rect 9824 16532 9830 16584
rect 9876 16572 9904 16603
rect 12434 16600 12440 16612
rect 12492 16600 12498 16652
rect 12544 16612 13216 16640
rect 11330 16572 11336 16584
rect 9876 16544 11336 16572
rect 11330 16532 11336 16544
rect 11388 16532 11394 16584
rect 12544 16581 12572 16612
rect 13188 16584 13216 16612
rect 13262 16600 13268 16652
rect 13320 16640 13326 16652
rect 15304 16649 15332 16736
rect 13357 16643 13415 16649
rect 13357 16640 13369 16643
rect 13320 16612 13369 16640
rect 13320 16600 13326 16612
rect 13357 16609 13369 16612
rect 13403 16609 13415 16643
rect 13357 16603 13415 16609
rect 15289 16643 15347 16649
rect 15289 16609 15301 16643
rect 15335 16609 15347 16643
rect 15289 16603 15347 16609
rect 15470 16600 15476 16652
rect 15528 16640 15534 16652
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 15528 16612 15761 16640
rect 15528 16600 15534 16612
rect 15749 16609 15761 16612
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 18322 16600 18328 16652
rect 18380 16640 18386 16652
rect 18601 16643 18659 16649
rect 18601 16640 18613 16643
rect 18380 16612 18613 16640
rect 18380 16600 18386 16612
rect 18601 16609 18613 16612
rect 18647 16640 18659 16643
rect 19242 16640 19248 16652
rect 18647 16612 19248 16640
rect 18647 16609 18659 16612
rect 18601 16603 18659 16609
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 19337 16643 19395 16649
rect 19337 16609 19349 16643
rect 19383 16640 19395 16643
rect 19797 16643 19855 16649
rect 19797 16640 19809 16643
rect 19383 16612 19809 16640
rect 19383 16609 19395 16612
rect 19337 16603 19395 16609
rect 19797 16609 19809 16612
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 20070 16600 20076 16652
rect 20128 16640 20134 16652
rect 20916 16649 20944 16736
rect 20349 16643 20407 16649
rect 20349 16640 20361 16643
rect 20128 16612 20361 16640
rect 20128 16600 20134 16612
rect 20349 16609 20361 16612
rect 20395 16609 20407 16643
rect 20901 16643 20959 16649
rect 20349 16603 20407 16609
rect 20456 16612 20760 16640
rect 12253 16575 12311 16581
rect 12253 16541 12265 16575
rect 12299 16572 12311 16575
rect 12529 16575 12587 16581
rect 12299 16544 12388 16572
rect 12299 16541 12311 16544
rect 12253 16535 12311 16541
rect 6871 16476 8248 16504
rect 6871 16473 6883 16476
rect 6825 16467 6883 16473
rect 1670 16396 1676 16448
rect 1728 16396 1734 16448
rect 3510 16396 3516 16448
rect 3568 16436 3574 16448
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 3568 16408 3801 16436
rect 3568 16396 3574 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 4798 16396 4804 16448
rect 4856 16396 4862 16448
rect 6748 16436 6776 16467
rect 8478 16464 8484 16516
rect 8536 16464 8542 16516
rect 9125 16507 9183 16513
rect 9125 16473 9137 16507
rect 9171 16473 9183 16507
rect 10106 16507 10164 16513
rect 10106 16504 10118 16507
rect 9125 16467 9183 16473
rect 9784 16476 10118 16504
rect 7466 16436 7472 16448
rect 6748 16408 7472 16436
rect 7466 16396 7472 16408
rect 7524 16396 7530 16448
rect 8570 16396 8576 16448
rect 8628 16436 8634 16448
rect 9140 16436 9168 16467
rect 9784 16445 9812 16476
rect 10106 16473 10118 16476
rect 10152 16473 10164 16507
rect 10106 16467 10164 16473
rect 12360 16448 12388 16544
rect 12529 16541 12541 16575
rect 12575 16541 12587 16575
rect 12529 16535 12587 16541
rect 12621 16575 12679 16581
rect 12621 16541 12633 16575
rect 12667 16572 12679 16575
rect 12710 16572 12716 16584
rect 12667 16544 12716 16572
rect 12667 16541 12679 16544
rect 12621 16535 12679 16541
rect 12710 16532 12716 16544
rect 12768 16572 12774 16584
rect 13081 16575 13139 16581
rect 13081 16572 13093 16575
rect 12768 16544 13093 16572
rect 12768 16532 12774 16544
rect 13081 16541 13093 16544
rect 13127 16541 13139 16575
rect 13081 16535 13139 16541
rect 12437 16507 12495 16513
rect 12437 16473 12449 16507
rect 12483 16473 12495 16507
rect 12437 16467 12495 16473
rect 8628 16408 9168 16436
rect 9769 16439 9827 16445
rect 8628 16396 8634 16408
rect 9769 16405 9781 16439
rect 9815 16405 9827 16439
rect 9769 16399 9827 16405
rect 11333 16439 11391 16445
rect 11333 16405 11345 16439
rect 11379 16436 11391 16439
rect 11422 16436 11428 16448
rect 11379 16408 11428 16436
rect 11379 16405 11391 16408
rect 11333 16399 11391 16405
rect 11422 16396 11428 16408
rect 11480 16396 11486 16448
rect 12342 16396 12348 16448
rect 12400 16396 12406 16448
rect 12452 16436 12480 16467
rect 12986 16464 12992 16516
rect 13044 16464 13050 16516
rect 13096 16504 13124 16535
rect 13170 16532 13176 16584
rect 13228 16532 13234 16584
rect 13446 16532 13452 16584
rect 13504 16572 13510 16584
rect 15488 16572 15516 16600
rect 13504 16544 15516 16572
rect 13504 16532 13510 16544
rect 15562 16532 15568 16584
rect 15620 16532 15626 16584
rect 17586 16532 17592 16584
rect 17644 16532 17650 16584
rect 17681 16575 17739 16581
rect 17681 16541 17693 16575
rect 17727 16541 17739 16575
rect 17681 16535 17739 16541
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16541 18935 16575
rect 18877 16535 18935 16541
rect 13354 16504 13360 16516
rect 13096 16476 13360 16504
rect 13354 16464 13360 16476
rect 13412 16464 13418 16516
rect 17696 16504 17724 16535
rect 18693 16507 18751 16513
rect 18693 16504 18705 16507
rect 17696 16476 18705 16504
rect 18693 16473 18705 16476
rect 18739 16473 18751 16507
rect 18892 16504 18920 16535
rect 19058 16532 19064 16584
rect 19116 16532 19122 16584
rect 19521 16575 19579 16581
rect 19521 16541 19533 16575
rect 19567 16572 19579 16575
rect 20456 16572 20484 16612
rect 20732 16581 20760 16612
rect 20901 16609 20913 16643
rect 20947 16609 20959 16643
rect 20901 16603 20959 16609
rect 19567 16544 20484 16572
rect 20717 16575 20775 16581
rect 19567 16541 19579 16544
rect 19521 16535 19579 16541
rect 19720 16504 19748 16544
rect 20717 16541 20729 16575
rect 20763 16541 20775 16575
rect 20717 16535 20775 16541
rect 21634 16532 21640 16584
rect 21692 16532 21698 16584
rect 18892 16476 19748 16504
rect 18693 16467 18751 16473
rect 12802 16436 12808 16448
rect 12452 16408 12808 16436
rect 12802 16396 12808 16408
rect 12860 16436 12866 16448
rect 13004 16436 13032 16464
rect 19720 16448 19748 16476
rect 12860 16408 13032 16436
rect 12860 16396 12866 16408
rect 14458 16396 14464 16448
rect 14516 16436 14522 16448
rect 14734 16436 14740 16448
rect 14516 16408 14740 16436
rect 14516 16396 14522 16408
rect 14734 16396 14740 16408
rect 14792 16436 14798 16448
rect 14829 16439 14887 16445
rect 14829 16436 14841 16439
rect 14792 16408 14841 16436
rect 14792 16396 14798 16408
rect 14829 16405 14841 16408
rect 14875 16405 14887 16439
rect 14829 16399 14887 16405
rect 17218 16396 17224 16448
rect 17276 16436 17282 16448
rect 17405 16439 17463 16445
rect 17405 16436 17417 16439
rect 17276 16408 17417 16436
rect 17276 16396 17282 16408
rect 17405 16405 17417 16408
rect 17451 16405 17463 16439
rect 17405 16399 17463 16405
rect 17957 16439 18015 16445
rect 17957 16405 17969 16439
rect 18003 16436 18015 16439
rect 18046 16436 18052 16448
rect 18003 16408 18052 16436
rect 18003 16405 18015 16408
rect 17957 16399 18015 16405
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 19702 16396 19708 16448
rect 19760 16396 19766 16448
rect 19978 16396 19984 16448
rect 20036 16436 20042 16448
rect 20533 16439 20591 16445
rect 20533 16436 20545 16439
rect 20036 16408 20545 16436
rect 20036 16396 20042 16408
rect 20533 16405 20545 16408
rect 20579 16405 20591 16439
rect 20533 16399 20591 16405
rect 20714 16396 20720 16448
rect 20772 16436 20778 16448
rect 20993 16439 21051 16445
rect 20993 16436 21005 16439
rect 20772 16408 21005 16436
rect 20772 16396 20778 16408
rect 20993 16405 21005 16408
rect 21039 16405 21051 16439
rect 20993 16399 21051 16405
rect 1104 16346 22264 16368
rect 1104 16294 4255 16346
rect 4307 16294 4319 16346
rect 4371 16294 4383 16346
rect 4435 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 9545 16346
rect 9597 16294 9609 16346
rect 9661 16294 9673 16346
rect 9725 16294 9737 16346
rect 9789 16294 9801 16346
rect 9853 16294 14835 16346
rect 14887 16294 14899 16346
rect 14951 16294 14963 16346
rect 15015 16294 15027 16346
rect 15079 16294 15091 16346
rect 15143 16294 20125 16346
rect 20177 16294 20189 16346
rect 20241 16294 20253 16346
rect 20305 16294 20317 16346
rect 20369 16294 20381 16346
rect 20433 16294 22264 16346
rect 1104 16272 22264 16294
rect 1670 16192 1676 16244
rect 1728 16232 1734 16244
rect 3053 16235 3111 16241
rect 3053 16232 3065 16235
rect 1728 16204 3065 16232
rect 1728 16192 1734 16204
rect 3053 16201 3065 16204
rect 3099 16232 3111 16235
rect 4614 16232 4620 16244
rect 3099 16204 4620 16232
rect 3099 16201 3111 16204
rect 3053 16195 3111 16201
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 5718 16192 5724 16244
rect 5776 16192 5782 16244
rect 6733 16235 6791 16241
rect 6733 16201 6745 16235
rect 6779 16232 6791 16235
rect 6914 16232 6920 16244
rect 6779 16204 6920 16232
rect 6779 16201 6791 16204
rect 6733 16195 6791 16201
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 9398 16232 9404 16244
rect 8352 16204 9404 16232
rect 8352 16192 8358 16204
rect 9398 16192 9404 16204
rect 9456 16192 9462 16244
rect 11790 16232 11796 16244
rect 9600 16204 11796 16232
rect 2130 16124 2136 16176
rect 2188 16164 2194 16176
rect 9600 16173 9628 16204
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 11977 16235 12035 16241
rect 11977 16201 11989 16235
rect 12023 16232 12035 16235
rect 14645 16235 14703 16241
rect 12023 16204 12357 16232
rect 12023 16201 12035 16204
rect 11977 16195 12035 16201
rect 2409 16167 2467 16173
rect 2409 16164 2421 16167
rect 2188 16136 2421 16164
rect 2188 16124 2194 16136
rect 2409 16133 2421 16136
rect 2455 16133 2467 16167
rect 2409 16127 2467 16133
rect 4341 16167 4399 16173
rect 4341 16133 4353 16167
rect 4387 16164 4399 16167
rect 9585 16167 9643 16173
rect 9585 16164 9597 16167
rect 4387 16136 9597 16164
rect 4387 16133 4399 16136
rect 4341 16127 4399 16133
rect 5368 16108 5396 16136
rect 9585 16133 9597 16136
rect 9631 16133 9643 16167
rect 9585 16127 9643 16133
rect 11088 16167 11146 16173
rect 11088 16133 11100 16167
rect 11134 16164 11146 16167
rect 11422 16164 11428 16176
rect 11134 16136 11428 16164
rect 11134 16133 11146 16136
rect 11088 16127 11146 16133
rect 11422 16124 11428 16136
rect 11480 16124 11486 16176
rect 11606 16124 11612 16176
rect 11664 16124 11670 16176
rect 12221 16167 12279 16173
rect 12221 16164 12233 16167
rect 11716 16136 12020 16164
rect 2314 16056 2320 16108
rect 2372 16056 2378 16108
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16096 2559 16099
rect 3234 16096 3240 16108
rect 2547 16068 3240 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 3234 16056 3240 16068
rect 3292 16056 3298 16108
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16065 4491 16099
rect 4433 16059 4491 16065
rect 4448 16028 4476 16059
rect 4522 16056 4528 16108
rect 4580 16096 4586 16108
rect 4617 16099 4675 16105
rect 4617 16096 4629 16099
rect 4580 16068 4629 16096
rect 4580 16056 4586 16068
rect 4617 16065 4629 16068
rect 4663 16065 4675 16099
rect 4617 16059 4675 16065
rect 4709 16099 4767 16105
rect 4709 16065 4721 16099
rect 4755 16065 4767 16099
rect 4709 16059 4767 16065
rect 4724 16028 4752 16059
rect 4798 16056 4804 16108
rect 4856 16056 4862 16108
rect 5258 16096 5264 16108
rect 4908 16068 5264 16096
rect 4908 16028 4936 16068
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 5350 16056 5356 16108
rect 5408 16056 5414 16108
rect 5905 16099 5963 16105
rect 5905 16065 5917 16099
rect 5951 16096 5963 16099
rect 6086 16096 6092 16108
rect 5951 16068 6092 16096
rect 5951 16065 5963 16068
rect 5905 16059 5963 16065
rect 6086 16056 6092 16068
rect 6144 16056 6150 16108
rect 6362 16056 6368 16108
rect 6420 16056 6426 16108
rect 6454 16056 6460 16108
rect 6512 16056 6518 16108
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 7098 16056 7104 16108
rect 7156 16096 7162 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 7156 16068 7389 16096
rect 7156 16056 7162 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 7466 16056 7472 16108
rect 7524 16056 7530 16108
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16065 7619 16099
rect 7561 16059 7619 16065
rect 4448 16000 4660 16028
rect 4724 16000 4936 16028
rect 5169 16031 5227 16037
rect 4632 15904 4660 16000
rect 5169 15997 5181 16031
rect 5215 16028 5227 16031
rect 5534 16028 5540 16040
rect 5215 16000 5540 16028
rect 5215 15997 5227 16000
rect 5169 15991 5227 15997
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 6181 16031 6239 16037
rect 6181 16028 6193 16031
rect 5644 16000 6193 16028
rect 4614 15852 4620 15904
rect 4672 15852 4678 15904
rect 4982 15852 4988 15904
rect 5040 15852 5046 15904
rect 5552 15892 5580 15988
rect 5644 15969 5672 16000
rect 6181 15997 6193 16000
rect 6227 16028 6239 16031
rect 6472 16028 6500 16056
rect 6227 16000 6500 16028
rect 7576 16028 7604 16059
rect 7650 16056 7656 16108
rect 7708 16096 7714 16108
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7708 16068 7757 16096
rect 7708 16056 7714 16068
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 7745 16059 7803 16065
rect 8202 16056 8208 16108
rect 8260 16056 8266 16108
rect 9214 16056 9220 16108
rect 9272 16096 9278 16108
rect 10318 16096 10324 16108
rect 9272 16068 10324 16096
rect 9272 16056 9278 16068
rect 10318 16056 10324 16068
rect 10376 16096 10382 16108
rect 10376 16068 11468 16096
rect 10376 16056 10382 16068
rect 8220 16028 8248 16056
rect 7576 16000 8248 16028
rect 6227 15997 6239 16000
rect 6181 15991 6239 15997
rect 11330 15988 11336 16040
rect 11388 15988 11394 16040
rect 11440 16028 11468 16068
rect 11514 16056 11520 16108
rect 11572 16096 11578 16108
rect 11716 16096 11744 16136
rect 11992 16118 12020 16136
rect 12155 16136 12233 16164
rect 12155 16118 12183 16136
rect 12221 16133 12233 16136
rect 12267 16133 12279 16167
rect 12221 16127 12279 16133
rect 11572 16068 11744 16096
rect 11793 16099 11851 16105
rect 11572 16056 11578 16068
rect 11793 16065 11805 16099
rect 11839 16065 11851 16099
rect 11992 16090 12183 16118
rect 11793 16059 11851 16065
rect 11808 16028 11836 16059
rect 11440 16000 11836 16028
rect 12329 16028 12357 16204
rect 14645 16201 14657 16235
rect 14691 16232 14703 16235
rect 15194 16232 15200 16244
rect 14691 16204 15200 16232
rect 14691 16201 14703 16204
rect 14645 16195 14703 16201
rect 15194 16192 15200 16204
rect 15252 16192 15258 16244
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 16209 16235 16267 16241
rect 16209 16232 16221 16235
rect 15528 16204 16221 16232
rect 15528 16192 15534 16204
rect 16209 16201 16221 16204
rect 16255 16201 16267 16235
rect 16209 16195 16267 16201
rect 19058 16192 19064 16244
rect 19116 16192 19122 16244
rect 19505 16235 19563 16241
rect 19505 16201 19517 16235
rect 19551 16232 19563 16235
rect 19794 16232 19800 16244
rect 19551 16204 19800 16232
rect 19551 16201 19563 16204
rect 19505 16195 19563 16201
rect 19794 16192 19800 16204
rect 19852 16192 19858 16244
rect 19978 16192 19984 16244
rect 20036 16192 20042 16244
rect 20165 16235 20223 16241
rect 20165 16201 20177 16235
rect 20211 16201 20223 16235
rect 20165 16195 20223 16201
rect 12437 16167 12495 16173
rect 12437 16133 12449 16167
rect 12483 16164 12495 16167
rect 12618 16164 12624 16176
rect 12483 16136 12624 16164
rect 12483 16133 12495 16136
rect 12437 16127 12495 16133
rect 12618 16124 12624 16136
rect 12676 16164 12682 16176
rect 14550 16164 14556 16176
rect 12676 16136 12940 16164
rect 12676 16124 12682 16136
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 12544 16028 12572 16059
rect 12710 16056 12716 16108
rect 12768 16056 12774 16108
rect 12802 16056 12808 16108
rect 12860 16056 12866 16108
rect 12912 16105 12940 16136
rect 14384 16136 14556 16164
rect 14384 16105 14412 16136
rect 14550 16124 14556 16136
rect 14608 16124 14614 16176
rect 19705 16167 19763 16173
rect 14844 16136 16988 16164
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16065 12955 16099
rect 14185 16099 14243 16105
rect 14185 16096 14197 16099
rect 12897 16059 12955 16065
rect 14016 16068 14197 16096
rect 12329 16000 12572 16028
rect 12989 16031 13047 16037
rect 5629 15963 5687 15969
rect 5629 15929 5641 15963
rect 5675 15929 5687 15963
rect 5629 15923 5687 15929
rect 6089 15963 6147 15969
rect 6089 15929 6101 15963
rect 6135 15960 6147 15963
rect 6638 15960 6644 15972
rect 6135 15932 6644 15960
rect 6135 15929 6147 15932
rect 6089 15923 6147 15929
rect 6638 15920 6644 15932
rect 6696 15960 6702 15972
rect 7101 15963 7159 15969
rect 7101 15960 7113 15963
rect 6696 15932 7113 15960
rect 6696 15920 6702 15932
rect 7101 15929 7113 15932
rect 7147 15929 7159 15963
rect 11808 15960 11836 16000
rect 12989 15997 13001 16031
rect 13035 16028 13047 16031
rect 13262 16028 13268 16040
rect 13035 16000 13268 16028
rect 13035 15997 13047 16000
rect 12989 15991 13047 15997
rect 13262 15988 13268 16000
rect 13320 15988 13326 16040
rect 11882 15960 11888 15972
rect 11808 15932 11888 15960
rect 7101 15923 7159 15929
rect 11882 15920 11888 15932
rect 11940 15920 11946 15972
rect 12066 15920 12072 15972
rect 12124 15920 12130 15972
rect 12434 15920 12440 15972
rect 12492 15960 12498 15972
rect 12529 15963 12587 15969
rect 12529 15960 12541 15963
rect 12492 15932 12541 15960
rect 12492 15920 12498 15932
rect 12529 15929 12541 15932
rect 12575 15929 12587 15963
rect 14016 15960 14044 16068
rect 14185 16065 14197 16068
rect 14231 16065 14243 16099
rect 14185 16059 14243 16065
rect 14369 16099 14427 16105
rect 14369 16065 14381 16099
rect 14415 16065 14427 16099
rect 14369 16059 14427 16065
rect 14458 16056 14464 16108
rect 14516 16056 14522 16108
rect 14642 16056 14648 16108
rect 14700 16096 14706 16108
rect 14737 16099 14795 16105
rect 14737 16096 14749 16099
rect 14700 16068 14749 16096
rect 14700 16056 14706 16068
rect 14737 16065 14749 16068
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 14090 15988 14096 16040
rect 14148 16028 14154 16040
rect 14844 16037 14872 16136
rect 16960 16108 16988 16136
rect 19705 16133 19717 16167
rect 19751 16133 19763 16167
rect 19705 16127 19763 16133
rect 14918 16056 14924 16108
rect 14976 16096 14982 16108
rect 15085 16099 15143 16105
rect 15085 16096 15097 16099
rect 14976 16068 15097 16096
rect 14976 16056 14982 16068
rect 15085 16065 15097 16068
rect 15131 16065 15143 16099
rect 15085 16059 15143 16065
rect 16942 16056 16948 16108
rect 17000 16056 17006 16108
rect 17218 16105 17224 16108
rect 17212 16096 17224 16105
rect 17179 16068 17224 16096
rect 17212 16059 17224 16068
rect 17218 16056 17224 16059
rect 17276 16056 17282 16108
rect 14829 16031 14887 16037
rect 14829 16028 14841 16031
rect 14148 16000 14841 16028
rect 14148 15988 14154 16000
rect 14829 15997 14841 16000
rect 14875 15997 14887 16031
rect 14829 15991 14887 15997
rect 18417 16031 18475 16037
rect 18417 15997 18429 16031
rect 18463 15997 18475 16031
rect 18417 15991 18475 15997
rect 14461 15963 14519 15969
rect 14461 15960 14473 15963
rect 14016 15932 14473 15960
rect 12529 15923 12587 15929
rect 14461 15929 14473 15932
rect 14507 15929 14519 15963
rect 14461 15923 14519 15929
rect 18432 15904 18460 15991
rect 19337 15963 19395 15969
rect 19337 15929 19349 15963
rect 19383 15960 19395 15963
rect 19610 15960 19616 15972
rect 19383 15932 19616 15960
rect 19383 15929 19395 15932
rect 19337 15923 19395 15929
rect 19610 15920 19616 15932
rect 19668 15920 19674 15972
rect 19720 15960 19748 16127
rect 19886 16056 19892 16108
rect 19944 16056 19950 16108
rect 19996 16105 20024 16192
rect 20180 16164 20208 16195
rect 20346 16192 20352 16244
rect 20404 16232 20410 16244
rect 21450 16232 21456 16244
rect 20404 16204 21456 16232
rect 20404 16192 20410 16204
rect 21450 16192 21456 16204
rect 21508 16192 21514 16244
rect 21634 16192 21640 16244
rect 21692 16192 21698 16244
rect 20502 16167 20560 16173
rect 20502 16164 20514 16167
rect 20180 16136 20514 16164
rect 20502 16133 20514 16136
rect 20548 16133 20560 16167
rect 20502 16127 20560 16133
rect 19981 16099 20039 16105
rect 19981 16065 19993 16099
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 19904 16028 19932 16056
rect 20257 16031 20315 16037
rect 20257 16028 20269 16031
rect 19904 16000 20269 16028
rect 20257 15997 20269 16000
rect 20303 15997 20315 16031
rect 20257 15991 20315 15997
rect 19720 15932 20300 15960
rect 20272 15904 20300 15932
rect 6546 15892 6552 15904
rect 5552 15864 6552 15892
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 9953 15895 10011 15901
rect 9953 15861 9965 15895
rect 9999 15892 10011 15895
rect 10134 15892 10140 15904
rect 9999 15864 10140 15892
rect 9999 15861 10011 15864
rect 9953 15855 10011 15861
rect 10134 15852 10140 15864
rect 10192 15892 10198 15904
rect 12250 15892 12256 15904
rect 10192 15864 12256 15892
rect 10192 15852 10198 15864
rect 12250 15852 12256 15864
rect 12308 15852 12314 15904
rect 14369 15895 14427 15901
rect 14369 15861 14381 15895
rect 14415 15892 14427 15895
rect 14826 15892 14832 15904
rect 14415 15864 14832 15892
rect 14415 15861 14427 15864
rect 14369 15855 14427 15861
rect 14826 15852 14832 15864
rect 14884 15852 14890 15904
rect 18325 15895 18383 15901
rect 18325 15861 18337 15895
rect 18371 15892 18383 15895
rect 18414 15892 18420 15904
rect 18371 15864 18420 15892
rect 18371 15861 18383 15864
rect 18325 15855 18383 15861
rect 18414 15852 18420 15864
rect 18472 15852 18478 15904
rect 19426 15852 19432 15904
rect 19484 15892 19490 15904
rect 19521 15895 19579 15901
rect 19521 15892 19533 15895
rect 19484 15864 19533 15892
rect 19484 15852 19490 15864
rect 19521 15861 19533 15864
rect 19567 15861 19579 15895
rect 19521 15855 19579 15861
rect 19702 15852 19708 15904
rect 19760 15892 19766 15904
rect 19886 15892 19892 15904
rect 19760 15864 19892 15892
rect 19760 15852 19766 15864
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 20254 15852 20260 15904
rect 20312 15852 20318 15904
rect 1104 15802 22264 15824
rect 1104 15750 3595 15802
rect 3647 15750 3659 15802
rect 3711 15750 3723 15802
rect 3775 15750 3787 15802
rect 3839 15750 3851 15802
rect 3903 15750 8885 15802
rect 8937 15750 8949 15802
rect 9001 15750 9013 15802
rect 9065 15750 9077 15802
rect 9129 15750 9141 15802
rect 9193 15750 14175 15802
rect 14227 15750 14239 15802
rect 14291 15750 14303 15802
rect 14355 15750 14367 15802
rect 14419 15750 14431 15802
rect 14483 15750 19465 15802
rect 19517 15750 19529 15802
rect 19581 15750 19593 15802
rect 19645 15750 19657 15802
rect 19709 15750 19721 15802
rect 19773 15750 22264 15802
rect 1104 15728 22264 15750
rect 2314 15648 2320 15700
rect 2372 15648 2378 15700
rect 3234 15688 3240 15700
rect 2424 15660 3240 15688
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15552 2283 15555
rect 2424 15552 2452 15660
rect 3234 15648 3240 15660
rect 3292 15648 3298 15700
rect 3510 15648 3516 15700
rect 3568 15648 3574 15700
rect 4525 15691 4583 15697
rect 4525 15657 4537 15691
rect 4571 15688 4583 15691
rect 4706 15688 4712 15700
rect 4571 15660 4712 15688
rect 4571 15657 4583 15660
rect 4525 15651 4583 15657
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 4982 15648 4988 15700
rect 5040 15648 5046 15700
rect 7282 15648 7288 15700
rect 7340 15688 7346 15700
rect 7469 15691 7527 15697
rect 7469 15688 7481 15691
rect 7340 15660 7481 15688
rect 7340 15648 7346 15660
rect 7469 15657 7481 15660
rect 7515 15657 7527 15691
rect 7469 15651 7527 15657
rect 7834 15648 7840 15700
rect 7892 15648 7898 15700
rect 11790 15648 11796 15700
rect 11848 15688 11854 15700
rect 12894 15688 12900 15700
rect 11848 15660 12900 15688
rect 11848 15648 11854 15660
rect 12894 15648 12900 15660
rect 12952 15648 12958 15700
rect 12989 15691 13047 15697
rect 12989 15657 13001 15691
rect 13035 15688 13047 15691
rect 13265 15691 13323 15697
rect 13265 15688 13277 15691
rect 13035 15660 13277 15688
rect 13035 15657 13047 15660
rect 12989 15651 13047 15657
rect 13265 15657 13277 15660
rect 13311 15657 13323 15691
rect 13265 15651 13323 15657
rect 14550 15648 14556 15700
rect 14608 15688 14614 15700
rect 14829 15691 14887 15697
rect 14829 15688 14841 15691
rect 14608 15660 14841 15688
rect 14608 15648 14614 15660
rect 14829 15657 14841 15660
rect 14875 15657 14887 15691
rect 14829 15651 14887 15657
rect 16942 15648 16948 15700
rect 17000 15648 17006 15700
rect 18141 15691 18199 15697
rect 18141 15657 18153 15691
rect 18187 15657 18199 15691
rect 18141 15651 18199 15657
rect 18785 15691 18843 15697
rect 18785 15657 18797 15691
rect 18831 15688 18843 15691
rect 19426 15688 19432 15700
rect 18831 15660 19432 15688
rect 18831 15657 18843 15660
rect 18785 15651 18843 15657
rect 3528 15620 3556 15648
rect 2271 15524 2452 15552
rect 2516 15592 3556 15620
rect 2271 15521 2283 15524
rect 2225 15515 2283 15521
rect 2516 15493 2544 15592
rect 3789 15555 3847 15561
rect 3789 15552 3801 15555
rect 2608 15524 3801 15552
rect 2608 15493 2636 15524
rect 3789 15521 3801 15524
rect 3835 15521 3847 15555
rect 3789 15515 3847 15521
rect 4062 15512 4068 15564
rect 4120 15552 4126 15564
rect 4522 15552 4528 15564
rect 4120 15524 4528 15552
rect 4120 15512 4126 15524
rect 4522 15512 4528 15524
rect 4580 15512 4586 15564
rect 5000 15552 5028 15648
rect 8570 15620 8576 15632
rect 4724 15524 5028 15552
rect 5276 15592 8576 15620
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15453 2467 15487
rect 2409 15447 2467 15453
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15453 2651 15487
rect 2593 15447 2651 15453
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15484 2743 15487
rect 3053 15487 3111 15493
rect 2731 15456 3004 15484
rect 2731 15453 2743 15456
rect 2685 15447 2743 15453
rect 2424 15416 2452 15447
rect 2700 15416 2728 15447
rect 2424 15388 2728 15416
rect 2869 15419 2927 15425
rect 2869 15385 2881 15419
rect 2915 15385 2927 15419
rect 2976 15416 3004 15456
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 4080 15484 4108 15512
rect 3099 15456 4108 15484
rect 4433 15487 4491 15493
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 4433 15453 4445 15487
rect 4479 15484 4491 15487
rect 4614 15484 4620 15496
rect 4479 15456 4620 15484
rect 4479 15453 4491 15456
rect 4433 15447 4491 15453
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 4724 15493 4752 15524
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15453 4767 15487
rect 4709 15447 4767 15453
rect 4982 15444 4988 15496
rect 5040 15444 5046 15496
rect 5276 15493 5304 15592
rect 8570 15580 8576 15592
rect 8628 15580 8634 15632
rect 13814 15620 13820 15632
rect 12912 15592 13820 15620
rect 8113 15555 8171 15561
rect 8113 15552 8125 15555
rect 7576 15524 8125 15552
rect 7576 15496 7604 15524
rect 8113 15521 8125 15524
rect 8159 15521 8171 15555
rect 8113 15515 8171 15521
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15552 8355 15555
rect 8386 15552 8392 15564
rect 8343 15524 8392 15552
rect 8343 15521 8355 15524
rect 8297 15515 8355 15521
rect 8386 15512 8392 15524
rect 8444 15552 8450 15564
rect 9214 15552 9220 15564
rect 8444 15524 9220 15552
rect 8444 15512 8450 15524
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 12342 15512 12348 15564
rect 12400 15552 12406 15564
rect 12912 15552 12940 15592
rect 13814 15580 13820 15592
rect 13872 15580 13878 15632
rect 18156 15620 18184 15651
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 19978 15648 19984 15700
rect 20036 15648 20042 15700
rect 20254 15648 20260 15700
rect 20312 15688 20318 15700
rect 21913 15691 21971 15697
rect 21913 15688 21925 15691
rect 20312 15660 21925 15688
rect 20312 15648 20318 15660
rect 21913 15657 21925 15660
rect 21959 15657 21971 15691
rect 21913 15651 21971 15657
rect 19886 15620 19892 15632
rect 18156 15592 19656 15620
rect 12400 15524 12940 15552
rect 12400 15512 12406 15524
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15453 5319 15487
rect 5261 15447 5319 15453
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 7558 15484 7564 15496
rect 7515 15456 7564 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 7650 15444 7656 15496
rect 7708 15444 7714 15496
rect 7745 15487 7803 15493
rect 7745 15453 7757 15487
rect 7791 15484 7803 15487
rect 8021 15487 8079 15493
rect 8021 15484 8033 15487
rect 7791 15456 8033 15484
rect 7791 15453 7803 15456
rect 7745 15447 7803 15453
rect 8021 15453 8033 15456
rect 8067 15453 8079 15487
rect 8021 15447 8079 15453
rect 8205 15487 8263 15493
rect 8205 15453 8217 15487
rect 8251 15453 8263 15487
rect 8205 15447 8263 15453
rect 3418 15416 3424 15428
rect 2976 15388 3424 15416
rect 2869 15379 2927 15385
rect 2590 15308 2596 15360
rect 2648 15308 2654 15360
rect 2884 15348 2912 15379
rect 3418 15376 3424 15388
rect 3476 15376 3482 15428
rect 5169 15419 5227 15425
rect 5169 15416 5181 15419
rect 4724 15388 5181 15416
rect 4724 15360 4752 15388
rect 5169 15385 5181 15388
rect 5215 15385 5227 15419
rect 7760 15416 7788 15447
rect 5169 15379 5227 15385
rect 7484 15388 7788 15416
rect 7484 15360 7512 15388
rect 3050 15348 3056 15360
rect 2884 15320 3056 15348
rect 3050 15308 3056 15320
rect 3108 15308 3114 15360
rect 3605 15351 3663 15357
rect 3605 15317 3617 15351
rect 3651 15348 3663 15351
rect 4154 15348 4160 15360
rect 3651 15320 4160 15348
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 4154 15308 4160 15320
rect 4212 15308 4218 15360
rect 4706 15308 4712 15360
rect 4764 15308 4770 15360
rect 4890 15308 4896 15360
rect 4948 15308 4954 15360
rect 7466 15308 7472 15360
rect 7524 15308 7530 15360
rect 7650 15308 7656 15360
rect 7708 15348 7714 15360
rect 8220 15348 8248 15447
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 12912 15484 12940 15524
rect 12986 15512 12992 15564
rect 13044 15552 13050 15564
rect 19628 15561 19656 15592
rect 19812 15592 19892 15620
rect 19613 15555 19671 15561
rect 13044 15524 15700 15552
rect 13044 15512 13050 15524
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 12216 15456 12848 15484
rect 12912 15456 13461 15484
rect 12216 15444 12222 15456
rect 12820 15416 12848 15456
rect 13449 15453 13461 15456
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15484 13691 15487
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 13679 15456 13737 15484
rect 13679 15453 13691 15456
rect 13633 15447 13691 15453
rect 13725 15453 13737 15456
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 13909 15487 13967 15493
rect 13909 15453 13921 15487
rect 13955 15484 13967 15487
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13955 15456 14105 15484
rect 13955 15453 13967 15456
rect 13909 15447 13967 15453
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 13173 15419 13231 15425
rect 13173 15416 13185 15419
rect 12820 15388 13185 15416
rect 13173 15385 13185 15388
rect 13219 15385 13231 15419
rect 13740 15416 13768 15447
rect 14274 15444 14280 15496
rect 14332 15484 14338 15496
rect 14645 15487 14703 15493
rect 14645 15484 14657 15487
rect 14332 15456 14657 15484
rect 14332 15444 14338 15456
rect 14645 15453 14657 15456
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 14826 15444 14832 15496
rect 14884 15484 14890 15496
rect 15013 15487 15071 15493
rect 15013 15484 15025 15487
rect 14884 15456 15025 15484
rect 14884 15444 14890 15456
rect 15013 15453 15025 15456
rect 15059 15453 15071 15487
rect 15013 15447 15071 15453
rect 15105 15487 15163 15493
rect 15105 15453 15117 15487
rect 15151 15453 15163 15487
rect 15105 15447 15163 15453
rect 13740 15388 13952 15416
rect 13173 15379 13231 15385
rect 7708 15320 8248 15348
rect 7708 15308 7714 15320
rect 12802 15308 12808 15360
rect 12860 15308 12866 15360
rect 12973 15351 13031 15357
rect 12973 15317 12985 15351
rect 13019 15348 13031 15351
rect 13078 15348 13084 15360
rect 13019 15320 13084 15348
rect 13019 15317 13031 15320
rect 12973 15311 13031 15317
rect 13078 15308 13084 15320
rect 13136 15348 13142 15360
rect 13817 15351 13875 15357
rect 13817 15348 13829 15351
rect 13136 15320 13829 15348
rect 13136 15308 13142 15320
rect 13817 15317 13829 15320
rect 13863 15317 13875 15351
rect 13924 15348 13952 15388
rect 14918 15376 14924 15428
rect 14976 15416 14982 15428
rect 15120 15416 15148 15447
rect 15194 15444 15200 15496
rect 15252 15444 15258 15496
rect 15286 15444 15292 15496
rect 15344 15444 15350 15496
rect 15672 15493 15700 15524
rect 19613 15521 19625 15555
rect 19659 15521 19671 15555
rect 19613 15515 19671 15521
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15453 15715 15487
rect 15657 15447 15715 15453
rect 16666 15444 16672 15496
rect 16724 15484 16730 15496
rect 17497 15487 17555 15493
rect 17497 15484 17509 15487
rect 16724 15456 17509 15484
rect 16724 15444 16730 15456
rect 17497 15453 17509 15456
rect 17543 15484 17555 15487
rect 18230 15484 18236 15496
rect 17543 15456 18236 15484
rect 17543 15453 17555 15456
rect 17497 15447 17555 15453
rect 18230 15444 18236 15456
rect 18288 15444 18294 15496
rect 18414 15444 18420 15496
rect 18472 15444 18478 15496
rect 19058 15444 19064 15496
rect 19116 15444 19122 15496
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15484 19487 15487
rect 19812 15484 19840 15592
rect 19886 15580 19892 15592
rect 19944 15580 19950 15632
rect 19996 15552 20024 15648
rect 20073 15555 20131 15561
rect 20073 15552 20085 15555
rect 19996 15524 20085 15552
rect 20073 15521 20085 15524
rect 20119 15521 20131 15555
rect 20073 15515 20131 15521
rect 19475 15456 19840 15484
rect 19475 15453 19487 15456
rect 19429 15447 19487 15453
rect 14976 15388 15148 15416
rect 14976 15376 14982 15388
rect 15212 15348 15240 15444
rect 15304 15416 15332 15444
rect 15746 15416 15752 15428
rect 15304 15388 15752 15416
rect 15746 15376 15752 15388
rect 15804 15376 15810 15428
rect 17586 15376 17592 15428
rect 17644 15416 17650 15428
rect 19245 15419 19303 15425
rect 19245 15416 19257 15419
rect 17644 15388 19257 15416
rect 17644 15376 17650 15388
rect 19245 15385 19257 15388
rect 19291 15385 19303 15419
rect 19444 15416 19472 15447
rect 19886 15444 19892 15496
rect 19944 15484 19950 15496
rect 19981 15487 20039 15493
rect 19981 15484 19993 15487
rect 19944 15456 19993 15484
rect 19944 15444 19950 15456
rect 19981 15453 19993 15456
rect 20027 15484 20039 15487
rect 20027 15456 20484 15484
rect 20027 15453 20039 15456
rect 19981 15447 20039 15453
rect 19610 15416 19616 15428
rect 19444 15388 19616 15416
rect 19245 15379 19303 15385
rect 19610 15376 19616 15388
rect 19668 15376 19674 15428
rect 19702 15376 19708 15428
rect 19760 15416 19766 15428
rect 20257 15419 20315 15425
rect 20257 15416 20269 15419
rect 19760 15388 20269 15416
rect 19760 15376 19766 15388
rect 20257 15385 20269 15388
rect 20303 15416 20315 15419
rect 20346 15416 20352 15428
rect 20303 15388 20352 15416
rect 20303 15385 20315 15388
rect 20257 15379 20315 15385
rect 20346 15376 20352 15388
rect 20404 15376 20410 15428
rect 20456 15416 20484 15456
rect 20530 15444 20536 15496
rect 20588 15444 20594 15496
rect 21634 15484 21640 15496
rect 20732 15456 21640 15484
rect 20732 15416 20760 15456
rect 21634 15444 21640 15456
rect 21692 15444 21698 15496
rect 20456 15388 20760 15416
rect 20800 15419 20858 15425
rect 20800 15385 20812 15419
rect 20846 15416 20858 15419
rect 20898 15416 20904 15428
rect 20846 15388 20904 15416
rect 20846 15385 20858 15388
rect 20800 15379 20858 15385
rect 20898 15376 20904 15388
rect 20956 15376 20962 15428
rect 13924 15320 15240 15348
rect 13817 15311 13875 15317
rect 18322 15308 18328 15360
rect 18380 15348 18386 15360
rect 18509 15351 18567 15357
rect 18509 15348 18521 15351
rect 18380 15320 18521 15348
rect 18380 15308 18386 15320
rect 18509 15317 18521 15320
rect 18555 15317 18567 15351
rect 18509 15311 18567 15317
rect 18598 15308 18604 15360
rect 18656 15308 18662 15360
rect 18874 15308 18880 15360
rect 18932 15308 18938 15360
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 19797 15351 19855 15357
rect 19797 15348 19809 15351
rect 19484 15320 19809 15348
rect 19484 15308 19490 15320
rect 19797 15317 19809 15320
rect 19843 15317 19855 15351
rect 19797 15311 19855 15317
rect 1104 15258 22264 15280
rect 1104 15206 4255 15258
rect 4307 15206 4319 15258
rect 4371 15206 4383 15258
rect 4435 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 9545 15258
rect 9597 15206 9609 15258
rect 9661 15206 9673 15258
rect 9725 15206 9737 15258
rect 9789 15206 9801 15258
rect 9853 15206 14835 15258
rect 14887 15206 14899 15258
rect 14951 15206 14963 15258
rect 15015 15206 15027 15258
rect 15079 15206 15091 15258
rect 15143 15206 20125 15258
rect 20177 15206 20189 15258
rect 20241 15206 20253 15258
rect 20305 15206 20317 15258
rect 20369 15206 20381 15258
rect 20433 15206 22264 15258
rect 1104 15184 22264 15206
rect 2777 15147 2835 15153
rect 2777 15113 2789 15147
rect 2823 15144 2835 15147
rect 2823 15116 4108 15144
rect 2823 15113 2835 15116
rect 2777 15107 2835 15113
rect 1664 15079 1722 15085
rect 1664 15045 1676 15079
rect 1710 15076 1722 15079
rect 2590 15076 2596 15088
rect 1710 15048 2596 15076
rect 1710 15045 1722 15048
rect 1664 15039 1722 15045
rect 2590 15036 2596 15048
rect 2648 15036 2654 15088
rect 3160 15085 3188 15116
rect 4080 15088 4108 15116
rect 4154 15104 4160 15156
rect 4212 15104 4218 15156
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 4982 15144 4988 15156
rect 4755 15116 4988 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 4982 15104 4988 15116
rect 5040 15104 5046 15156
rect 12802 15144 12808 15156
rect 12176 15116 12808 15144
rect 3145 15079 3203 15085
rect 3145 15045 3157 15079
rect 3191 15045 3203 15079
rect 3145 15039 3203 15045
rect 3361 15079 3419 15085
rect 3361 15045 3373 15079
rect 3407 15076 3419 15079
rect 3510 15076 3516 15088
rect 3407 15048 3516 15076
rect 3407 15045 3419 15048
rect 3361 15039 3419 15045
rect 3510 15036 3516 15048
rect 3568 15036 3574 15088
rect 4062 15036 4068 15088
rect 4120 15036 4126 15088
rect 4172 15076 4200 15104
rect 4801 15079 4859 15085
rect 4801 15076 4813 15079
rect 4172 15048 4813 15076
rect 4801 15045 4813 15048
rect 4847 15045 4859 15079
rect 4801 15039 4859 15045
rect 6457 15079 6515 15085
rect 6457 15045 6469 15079
rect 6503 15076 6515 15079
rect 6546 15076 6552 15088
rect 6503 15048 6552 15076
rect 6503 15045 6515 15048
rect 6457 15039 6515 15045
rect 6546 15036 6552 15048
rect 6604 15076 6610 15088
rect 8478 15076 8484 15088
rect 6604 15048 8484 15076
rect 6604 15036 6610 15048
rect 8478 15036 8484 15048
rect 8536 15036 8542 15088
rect 1397 15011 1455 15017
rect 1397 14977 1409 15011
rect 1443 15008 1455 15011
rect 1486 15008 1492 15020
rect 1443 14980 1492 15008
rect 1443 14977 1455 14980
rect 1397 14971 1455 14977
rect 1486 14968 1492 14980
rect 1544 14968 1550 15020
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 14977 3847 15011
rect 3789 14971 3847 14977
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 15008 4215 15011
rect 4203 14980 4384 15008
rect 4203 14977 4215 14980
rect 4157 14971 4215 14977
rect 3142 14900 3148 14952
rect 3200 14940 3206 14952
rect 3605 14943 3663 14949
rect 3605 14940 3617 14943
rect 3200 14912 3617 14940
rect 3200 14900 3206 14912
rect 3605 14909 3617 14912
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 3418 14832 3424 14884
rect 3476 14872 3482 14884
rect 3513 14875 3571 14881
rect 3513 14872 3525 14875
rect 3476 14844 3525 14872
rect 3476 14832 3482 14844
rect 3513 14841 3525 14844
rect 3559 14841 3571 14875
rect 3804 14872 3832 14971
rect 4062 14900 4068 14952
rect 4120 14900 4126 14952
rect 4246 14900 4252 14952
rect 4304 14900 4310 14952
rect 4356 14940 4384 14980
rect 4430 14968 4436 15020
rect 4488 14968 4494 15020
rect 4522 14968 4528 15020
rect 4580 15008 4586 15020
rect 4985 15011 5043 15017
rect 4985 15008 4997 15011
rect 4580 14980 4997 15008
rect 4580 14968 4586 14980
rect 4985 14977 4997 14980
rect 5031 14977 5043 15011
rect 4985 14971 5043 14977
rect 5077 15011 5135 15017
rect 5077 14977 5089 15011
rect 5123 14977 5135 15011
rect 5077 14971 5135 14977
rect 4356 14912 4476 14940
rect 4448 14872 4476 14912
rect 4614 14900 4620 14952
rect 4672 14940 4678 14952
rect 4672 14912 4844 14940
rect 4672 14900 4678 14912
rect 4706 14872 4712 14884
rect 3804 14844 4108 14872
rect 4448 14844 4712 14872
rect 3513 14835 3571 14841
rect 3326 14764 3332 14816
rect 3384 14764 3390 14816
rect 3970 14764 3976 14816
rect 4028 14764 4034 14816
rect 4080 14804 4108 14844
rect 4706 14832 4712 14844
rect 4764 14832 4770 14884
rect 4816 14881 4844 14912
rect 4801 14875 4859 14881
rect 4801 14841 4813 14875
rect 4847 14841 4859 14875
rect 4801 14835 4859 14841
rect 5092 14816 5120 14971
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 8386 15008 8392 15020
rect 6788 14980 8392 15008
rect 6788 14968 6794 14980
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 12176 15017 12204 15116
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 14274 15144 14280 15156
rect 13872 15116 14280 15144
rect 13872 15104 13878 15116
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 14642 15104 14648 15156
rect 14700 15144 14706 15156
rect 14737 15147 14795 15153
rect 14737 15144 14749 15147
rect 14700 15116 14749 15144
rect 14700 15104 14706 15116
rect 14737 15113 14749 15116
rect 14783 15113 14795 15147
rect 14737 15107 14795 15113
rect 15473 15147 15531 15153
rect 15473 15113 15485 15147
rect 15519 15144 15531 15147
rect 15562 15144 15568 15156
rect 15519 15116 15568 15144
rect 15519 15113 15531 15116
rect 15473 15107 15531 15113
rect 15562 15104 15568 15116
rect 15620 15104 15626 15156
rect 16666 15104 16672 15156
rect 16724 15104 16730 15156
rect 18874 15144 18880 15156
rect 18156 15116 18880 15144
rect 14090 15076 14096 15088
rect 12452 15048 14096 15076
rect 12452 15017 12480 15048
rect 14090 15036 14096 15048
rect 14148 15036 14154 15088
rect 14292 15017 14320 15104
rect 16960 15048 18092 15076
rect 16960 15020 16988 15048
rect 12161 15011 12219 15017
rect 12161 14977 12173 15011
rect 12207 14977 12219 15011
rect 12161 14971 12219 14977
rect 12437 15011 12495 15017
rect 12437 14977 12449 15011
rect 12483 14977 12495 15011
rect 12693 15011 12751 15017
rect 12693 15008 12705 15011
rect 12437 14971 12495 14977
rect 12544 14980 12705 15008
rect 12544 14940 12572 14980
rect 12693 14977 12705 14980
rect 12739 14977 12751 15011
rect 12693 14971 12751 14977
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 15008 14611 15011
rect 15194 15008 15200 15020
rect 14599 14980 15200 15008
rect 14599 14977 14611 14980
rect 14553 14971 14611 14977
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 15562 14968 15568 15020
rect 15620 14968 15626 15020
rect 16942 14968 16948 15020
rect 17000 14968 17006 15020
rect 18064 15017 18092 15048
rect 17793 15011 17851 15017
rect 17793 14977 17805 15011
rect 17839 15008 17851 15011
rect 18049 15011 18107 15017
rect 17839 14980 18000 15008
rect 17839 14977 17851 14980
rect 17793 14971 17851 14977
rect 12360 14912 12572 14940
rect 17972 14940 18000 14980
rect 18049 14977 18061 15011
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 18156 14940 18184 15116
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 19702 15104 19708 15156
rect 19760 15104 19766 15156
rect 19794 15104 19800 15156
rect 19852 15104 19858 15156
rect 20714 15144 20720 15156
rect 20272 15116 20720 15144
rect 18233 15079 18291 15085
rect 18233 15045 18245 15079
rect 18279 15076 18291 15079
rect 18598 15076 18604 15088
rect 18279 15048 18604 15076
rect 18279 15045 18291 15048
rect 18233 15039 18291 15045
rect 18598 15036 18604 15048
rect 18656 15036 18662 15088
rect 19334 15076 19340 15088
rect 18800 15048 19340 15076
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 18800 15017 18828 15048
rect 19334 15036 19340 15048
rect 19392 15036 19398 15088
rect 19720 15076 19748 15104
rect 19949 15079 20007 15085
rect 19949 15076 19961 15079
rect 19720 15048 19961 15076
rect 19949 15045 19961 15048
rect 19995 15045 20007 15079
rect 19949 15039 20007 15045
rect 20165 15079 20223 15085
rect 20165 15045 20177 15079
rect 20211 15045 20223 15079
rect 20165 15039 20223 15045
rect 18417 15011 18475 15017
rect 18417 15008 18429 15011
rect 18380 14980 18429 15008
rect 18380 14968 18386 14980
rect 18417 14977 18429 14980
rect 18463 14977 18475 15011
rect 18417 14971 18475 14977
rect 18509 15011 18567 15017
rect 18509 14977 18521 15011
rect 18555 14977 18567 15011
rect 18509 14971 18567 14977
rect 18785 15011 18843 15017
rect 18785 14977 18797 15011
rect 18831 14977 18843 15011
rect 18785 14971 18843 14977
rect 19061 15011 19119 15017
rect 19061 14977 19073 15011
rect 19107 14977 19119 15011
rect 19061 14971 19119 14977
rect 19245 15011 19303 15017
rect 19245 14977 19257 15011
rect 19291 15008 19303 15011
rect 19426 15008 19432 15020
rect 19291 14980 19432 15008
rect 19291 14977 19303 14980
rect 19245 14971 19303 14977
rect 17972 14912 18184 14940
rect 7006 14832 7012 14884
rect 7064 14872 7070 14884
rect 7650 14872 7656 14884
rect 7064 14844 7656 14872
rect 7064 14832 7070 14844
rect 7650 14832 7656 14844
rect 7708 14832 7714 14884
rect 12360 14881 12388 14912
rect 18230 14900 18236 14952
rect 18288 14940 18294 14952
rect 18524 14940 18552 14971
rect 19076 14940 19104 14971
rect 19426 14968 19432 14980
rect 19484 14968 19490 15020
rect 19521 15011 19579 15017
rect 19521 14977 19533 15011
rect 19567 14977 19579 15011
rect 19521 14971 19579 14977
rect 18288 14912 18552 14940
rect 18708 14912 19104 14940
rect 18288 14900 18294 14912
rect 18708 14881 18736 14912
rect 12345 14875 12403 14881
rect 12345 14841 12357 14875
rect 12391 14841 12403 14875
rect 12345 14835 12403 14841
rect 18693 14875 18751 14881
rect 18693 14841 18705 14875
rect 18739 14841 18751 14875
rect 18693 14835 18751 14841
rect 18969 14875 19027 14881
rect 18969 14841 18981 14875
rect 19015 14872 19027 14875
rect 19242 14872 19248 14884
rect 19015 14844 19248 14872
rect 19015 14841 19027 14844
rect 18969 14835 19027 14841
rect 19242 14832 19248 14844
rect 19300 14872 19306 14884
rect 19536 14872 19564 14971
rect 19886 14900 19892 14952
rect 19944 14940 19950 14952
rect 20180 14940 20208 15039
rect 20272 15017 20300 15116
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 20898 15104 20904 15156
rect 20956 15104 20962 15156
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 20441 15011 20499 15017
rect 20441 14977 20453 15011
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 20625 15011 20683 15017
rect 20625 14977 20637 15011
rect 20671 15008 20683 15011
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 20671 14980 20729 15008
rect 20671 14977 20683 14980
rect 20625 14971 20683 14977
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 19944 14912 20208 14940
rect 19944 14900 19950 14912
rect 19300 14844 19564 14872
rect 19300 14832 19306 14844
rect 19610 14832 19616 14884
rect 19668 14872 19674 14884
rect 20456 14872 20484 14971
rect 19668 14844 20484 14872
rect 19668 14832 19674 14844
rect 19904 14816 19932 14844
rect 4154 14804 4160 14816
rect 4080 14776 4160 14804
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 5074 14764 5080 14816
rect 5132 14764 5138 14816
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 6733 14807 6791 14813
rect 6733 14804 6745 14807
rect 5868 14776 6745 14804
rect 5868 14764 5874 14776
rect 6733 14773 6745 14776
rect 6779 14804 6791 14807
rect 6822 14804 6828 14816
rect 6779 14776 6828 14804
rect 6779 14773 6791 14776
rect 6733 14767 6791 14773
rect 6822 14764 6828 14776
rect 6880 14804 6886 14816
rect 7374 14804 7380 14816
rect 6880 14776 7380 14804
rect 6880 14764 6886 14776
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 14369 14807 14427 14813
rect 14369 14773 14381 14807
rect 14415 14804 14427 14807
rect 14550 14804 14556 14816
rect 14415 14776 14556 14804
rect 14415 14773 14427 14776
rect 14369 14767 14427 14773
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 18414 14764 18420 14816
rect 18472 14764 18478 14816
rect 19334 14764 19340 14816
rect 19392 14804 19398 14816
rect 19705 14807 19763 14813
rect 19705 14804 19717 14807
rect 19392 14776 19717 14804
rect 19392 14764 19398 14776
rect 19705 14773 19717 14776
rect 19751 14773 19763 14807
rect 19705 14767 19763 14773
rect 19886 14764 19892 14816
rect 19944 14764 19950 14816
rect 19978 14764 19984 14816
rect 20036 14764 20042 14816
rect 1104 14714 22264 14736
rect 1104 14662 3595 14714
rect 3647 14662 3659 14714
rect 3711 14662 3723 14714
rect 3775 14662 3787 14714
rect 3839 14662 3851 14714
rect 3903 14662 8885 14714
rect 8937 14662 8949 14714
rect 9001 14662 9013 14714
rect 9065 14662 9077 14714
rect 9129 14662 9141 14714
rect 9193 14662 14175 14714
rect 14227 14662 14239 14714
rect 14291 14662 14303 14714
rect 14355 14662 14367 14714
rect 14419 14662 14431 14714
rect 14483 14662 19465 14714
rect 19517 14662 19529 14714
rect 19581 14662 19593 14714
rect 19645 14662 19657 14714
rect 19709 14662 19721 14714
rect 19773 14662 22264 14714
rect 1104 14640 22264 14662
rect 3142 14560 3148 14612
rect 3200 14560 3206 14612
rect 3326 14560 3332 14612
rect 3384 14600 3390 14612
rect 3421 14603 3479 14609
rect 3421 14600 3433 14603
rect 3384 14572 3433 14600
rect 3384 14560 3390 14572
rect 3421 14569 3433 14572
rect 3467 14569 3479 14603
rect 3421 14563 3479 14569
rect 3881 14603 3939 14609
rect 3881 14569 3893 14603
rect 3927 14600 3939 14603
rect 4062 14600 4068 14612
rect 3927 14572 4068 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 1486 14424 1492 14476
rect 1544 14464 1550 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1544 14436 2053 14464
rect 1544 14424 1550 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 2308 14399 2366 14405
rect 2308 14365 2320 14399
rect 2354 14396 2366 14399
rect 3160 14396 3188 14560
rect 3436 14464 3464 14563
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 4430 14560 4436 14612
rect 4488 14560 4494 14612
rect 4890 14560 4896 14612
rect 4948 14600 4954 14612
rect 5353 14603 5411 14609
rect 5353 14600 5365 14603
rect 4948 14572 5365 14600
rect 4948 14560 4954 14572
rect 5353 14569 5365 14572
rect 5399 14569 5411 14603
rect 5353 14563 5411 14569
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 7837 14603 7895 14609
rect 7837 14600 7849 14603
rect 7524 14572 7849 14600
rect 7524 14560 7530 14572
rect 7837 14569 7849 14572
rect 7883 14569 7895 14603
rect 7837 14563 7895 14569
rect 8478 14560 8484 14612
rect 8536 14600 8542 14612
rect 9677 14603 9735 14609
rect 9677 14600 9689 14603
rect 8536 14572 9689 14600
rect 8536 14560 8542 14572
rect 9677 14569 9689 14572
rect 9723 14569 9735 14603
rect 9677 14563 9735 14569
rect 12989 14603 13047 14609
rect 12989 14569 13001 14603
rect 13035 14600 13047 14603
rect 13035 14572 13492 14600
rect 13035 14569 13047 14572
rect 12989 14563 13047 14569
rect 4448 14532 4476 14560
rect 4448 14504 5672 14532
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 3436 14436 4445 14464
rect 4433 14433 4445 14436
rect 4479 14464 4491 14467
rect 4522 14464 4528 14476
rect 4479 14436 4528 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4522 14424 4528 14436
rect 4580 14464 4586 14476
rect 5442 14464 5448 14476
rect 4580 14436 5448 14464
rect 4580 14424 4586 14436
rect 5442 14424 5448 14436
rect 5500 14464 5506 14476
rect 5644 14464 5672 14504
rect 5994 14492 6000 14544
rect 6052 14492 6058 14544
rect 8662 14532 8668 14544
rect 6104 14504 8668 14532
rect 6104 14464 6132 14504
rect 8662 14492 8668 14504
rect 8720 14492 8726 14544
rect 8754 14492 8760 14544
rect 8812 14532 8818 14544
rect 9125 14535 9183 14541
rect 8812 14504 9076 14532
rect 8812 14492 8818 14504
rect 7834 14464 7840 14476
rect 5500 14436 5580 14464
rect 5500 14424 5506 14436
rect 2354 14368 3188 14396
rect 2354 14365 2366 14368
rect 2308 14359 2366 14365
rect 3510 14356 3516 14408
rect 3568 14396 3574 14408
rect 5074 14396 5080 14408
rect 3568 14368 5080 14396
rect 3568 14356 3574 14368
rect 5074 14356 5080 14368
rect 5132 14396 5138 14408
rect 5552 14405 5580 14436
rect 5644 14436 6132 14464
rect 6196 14436 7236 14464
rect 5644 14408 5672 14436
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 5132 14368 5181 14396
rect 5132 14356 5138 14368
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 5537 14399 5595 14405
rect 5537 14365 5549 14399
rect 5583 14365 5595 14399
rect 5537 14359 5595 14365
rect 3970 14288 3976 14340
rect 4028 14328 4034 14340
rect 4617 14331 4675 14337
rect 4617 14328 4629 14331
rect 4028 14300 4629 14328
rect 4028 14288 4034 14300
rect 4617 14297 4629 14300
rect 4663 14297 4675 14331
rect 5184 14328 5212 14359
rect 5626 14356 5632 14408
rect 5684 14356 5690 14408
rect 6196 14405 6224 14436
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 5905 14399 5963 14405
rect 5905 14365 5917 14399
rect 5951 14396 5963 14399
rect 6181 14399 6239 14405
rect 6181 14396 6193 14399
rect 5951 14368 6193 14396
rect 5951 14365 5963 14368
rect 5905 14359 5963 14365
rect 6181 14365 6193 14368
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 6273 14399 6331 14405
rect 6273 14365 6285 14399
rect 6319 14396 6331 14399
rect 6319 14368 6684 14396
rect 6319 14365 6331 14368
rect 6273 14359 6331 14365
rect 5828 14328 5856 14359
rect 5184 14300 5856 14328
rect 5997 14331 6055 14337
rect 4617 14291 4675 14297
rect 5997 14297 6009 14331
rect 6043 14328 6055 14331
rect 6549 14331 6607 14337
rect 6549 14328 6561 14331
rect 6043 14300 6561 14328
rect 6043 14297 6055 14300
rect 5997 14291 6055 14297
rect 6549 14297 6561 14300
rect 6595 14297 6607 14331
rect 6549 14291 6607 14297
rect 6656 14260 6684 14368
rect 6730 14356 6736 14408
rect 6788 14356 6794 14408
rect 7006 14356 7012 14408
rect 7064 14356 7070 14408
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14365 7159 14399
rect 7101 14359 7159 14365
rect 6914 14288 6920 14340
rect 6972 14328 6978 14340
rect 7116 14328 7144 14359
rect 7208 14337 7236 14436
rect 7668 14436 7840 14464
rect 7466 14356 7472 14408
rect 7524 14356 7530 14408
rect 7668 14405 7696 14436
rect 7834 14424 7840 14436
rect 7892 14464 7898 14476
rect 8941 14467 8999 14473
rect 8941 14464 8953 14467
rect 7892 14436 8953 14464
rect 7892 14424 7898 14436
rect 8941 14433 8953 14436
rect 8987 14433 8999 14467
rect 9048 14464 9076 14504
rect 9125 14501 9137 14535
rect 9171 14532 9183 14535
rect 9214 14532 9220 14544
rect 9171 14504 9220 14532
rect 9171 14501 9183 14504
rect 9125 14495 9183 14501
rect 9214 14492 9220 14504
rect 9272 14492 9278 14544
rect 13173 14535 13231 14541
rect 13173 14501 13185 14535
rect 13219 14501 13231 14535
rect 13173 14495 13231 14501
rect 13188 14464 13216 14495
rect 9048 14436 9674 14464
rect 8941 14427 8999 14433
rect 7653 14399 7711 14405
rect 7653 14365 7665 14399
rect 7699 14365 7711 14399
rect 7653 14359 7711 14365
rect 8018 14356 8024 14408
rect 8076 14356 8082 14408
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 8386 14396 8392 14408
rect 8343 14368 8392 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 8481 14399 8539 14405
rect 8481 14365 8493 14399
rect 8527 14396 8539 14399
rect 8573 14399 8631 14405
rect 8573 14396 8585 14399
rect 8527 14368 8585 14396
rect 8527 14365 8539 14368
rect 8481 14359 8539 14365
rect 8573 14365 8585 14368
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 6972 14300 7144 14328
rect 7193 14331 7251 14337
rect 6972 14288 6978 14300
rect 7193 14297 7205 14331
rect 7239 14328 7251 14331
rect 7239 14300 8432 14328
rect 7239 14297 7251 14300
rect 7193 14291 7251 14297
rect 8404 14272 8432 14300
rect 8496 14272 8524 14359
rect 9490 14356 9496 14408
rect 9548 14356 9554 14408
rect 9306 14288 9312 14340
rect 9364 14328 9370 14340
rect 9401 14331 9459 14337
rect 9401 14328 9413 14331
rect 9364 14300 9413 14328
rect 9364 14288 9370 14300
rect 9401 14297 9413 14300
rect 9447 14297 9459 14331
rect 9646 14328 9674 14436
rect 9876 14436 10272 14464
rect 9876 14405 9904 14436
rect 10244 14408 10272 14436
rect 12820 14436 13216 14464
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14365 9919 14399
rect 9861 14359 9919 14365
rect 10045 14399 10103 14405
rect 10045 14365 10057 14399
rect 10091 14396 10103 14399
rect 10134 14396 10140 14408
rect 10091 14368 10140 14396
rect 10091 14365 10103 14368
rect 10045 14359 10103 14365
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 10226 14356 10232 14408
rect 10284 14356 10290 14408
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14396 10747 14399
rect 10962 14396 10968 14408
rect 10735 14368 10968 14396
rect 10735 14365 10747 14368
rect 10689 14359 10747 14365
rect 10962 14356 10968 14368
rect 11020 14356 11026 14408
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14396 11207 14399
rect 11882 14396 11888 14408
rect 11195 14368 11888 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11882 14356 11888 14368
rect 11940 14396 11946 14408
rect 12158 14396 12164 14408
rect 11940 14368 12164 14396
rect 11940 14356 11946 14368
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 12820 14405 12848 14436
rect 12805 14399 12863 14405
rect 12805 14365 12817 14399
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13464 14405 13492 14572
rect 14550 14560 14556 14612
rect 14608 14560 14614 14612
rect 14737 14603 14795 14609
rect 14737 14569 14749 14603
rect 14783 14569 14795 14603
rect 14737 14563 14795 14569
rect 13722 14424 13728 14476
rect 13780 14464 13786 14476
rect 14752 14464 14780 14563
rect 15194 14560 15200 14612
rect 15252 14560 15258 14612
rect 18046 14600 18052 14612
rect 16592 14572 18052 14600
rect 16298 14532 16304 14544
rect 15580 14504 16304 14532
rect 15286 14464 15292 14476
rect 13780 14436 14504 14464
rect 14752 14436 15292 14464
rect 13780 14424 13786 14436
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 13136 14368 13369 14396
rect 13136 14356 13142 14368
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 13449 14399 13507 14405
rect 13449 14365 13461 14399
rect 13495 14396 13507 14399
rect 13495 14368 14412 14396
rect 13495 14365 13507 14368
rect 13449 14359 13507 14365
rect 13173 14331 13231 14337
rect 13173 14328 13185 14331
rect 9646 14300 13185 14328
rect 9401 14291 9459 14297
rect 13173 14297 13185 14300
rect 13219 14297 13231 14331
rect 13173 14291 13231 14297
rect 14384 14272 14412 14368
rect 14476 14328 14504 14436
rect 15286 14424 15292 14436
rect 15344 14464 15350 14476
rect 15381 14467 15439 14473
rect 15381 14464 15393 14467
rect 15344 14436 15393 14464
rect 15344 14424 15350 14436
rect 15381 14433 15393 14436
rect 15427 14433 15439 14467
rect 15381 14427 15439 14433
rect 14642 14356 14648 14408
rect 14700 14396 14706 14408
rect 15105 14399 15163 14405
rect 15105 14396 15117 14399
rect 14700 14368 15117 14396
rect 14700 14356 14706 14368
rect 15105 14365 15117 14368
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 15470 14356 15476 14408
rect 15528 14356 15534 14408
rect 15580 14405 15608 14504
rect 16298 14492 16304 14504
rect 16356 14492 16362 14544
rect 16592 14473 16620 14572
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 18417 14603 18475 14609
rect 18417 14569 18429 14603
rect 18463 14600 18475 14603
rect 18598 14600 18604 14612
rect 18463 14572 18604 14600
rect 18463 14569 18475 14572
rect 18417 14563 18475 14569
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 19242 14600 19248 14612
rect 19168 14572 19248 14600
rect 15657 14467 15715 14473
rect 15657 14433 15669 14467
rect 15703 14433 15715 14467
rect 15657 14427 15715 14433
rect 16577 14467 16635 14473
rect 16577 14433 16589 14467
rect 16623 14433 16635 14467
rect 16577 14427 16635 14433
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 14737 14331 14795 14337
rect 14737 14328 14749 14331
rect 14476 14300 14749 14328
rect 14737 14297 14749 14300
rect 14783 14328 14795 14331
rect 15672 14328 15700 14427
rect 16942 14424 16948 14476
rect 17000 14464 17006 14476
rect 17037 14467 17095 14473
rect 17037 14464 17049 14467
rect 17000 14436 17049 14464
rect 17000 14424 17006 14436
rect 17037 14433 17049 14436
rect 17083 14433 17095 14467
rect 17037 14427 17095 14433
rect 16758 14356 16764 14408
rect 16816 14356 16822 14408
rect 19168 14396 19196 14572
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19334 14560 19340 14612
rect 19392 14560 19398 14612
rect 19352 14532 19380 14560
rect 19260 14504 19380 14532
rect 19260 14473 19288 14504
rect 19245 14467 19303 14473
rect 19245 14433 19257 14467
rect 19291 14433 19303 14467
rect 19245 14427 19303 14433
rect 19521 14399 19579 14405
rect 19521 14396 19533 14399
rect 19168 14368 19533 14396
rect 19521 14365 19533 14368
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 17304 14331 17362 14337
rect 14783 14300 15700 14328
rect 16040 14300 17080 14328
rect 14783 14297 14795 14300
rect 14737 14291 14795 14297
rect 7469 14263 7527 14269
rect 7469 14260 7481 14263
rect 6656 14232 7481 14260
rect 7469 14229 7481 14232
rect 7515 14260 7527 14263
rect 7742 14260 7748 14272
rect 7515 14232 7748 14260
rect 7515 14229 7527 14232
rect 7469 14223 7527 14229
rect 7742 14220 7748 14232
rect 7800 14220 7806 14272
rect 8386 14220 8392 14272
rect 8444 14220 8450 14272
rect 8478 14220 8484 14272
rect 8536 14220 8542 14272
rect 9953 14263 10011 14269
rect 9953 14229 9965 14263
rect 9999 14260 10011 14263
rect 10042 14260 10048 14272
rect 9999 14232 10048 14260
rect 9999 14229 10011 14232
rect 9953 14223 10011 14229
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 10870 14220 10876 14272
rect 10928 14220 10934 14272
rect 11333 14263 11391 14269
rect 11333 14229 11345 14263
rect 11379 14260 11391 14263
rect 11606 14260 11612 14272
rect 11379 14232 11612 14260
rect 11379 14229 11391 14232
rect 11333 14223 11391 14229
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 12618 14220 12624 14272
rect 12676 14220 12682 14272
rect 14366 14220 14372 14272
rect 14424 14220 14430 14272
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 16040 14260 16068 14300
rect 14516 14232 16068 14260
rect 14516 14220 14522 14232
rect 16942 14220 16948 14272
rect 17000 14220 17006 14272
rect 17052 14260 17080 14300
rect 17304 14297 17316 14331
rect 17350 14328 17362 14331
rect 17586 14328 17592 14340
rect 17350 14300 17592 14328
rect 17350 14297 17362 14300
rect 17304 14291 17362 14297
rect 17586 14288 17592 14300
rect 17644 14288 17650 14340
rect 20257 14263 20315 14269
rect 20257 14260 20269 14263
rect 17052 14232 20269 14260
rect 20257 14229 20269 14232
rect 20303 14229 20315 14263
rect 20257 14223 20315 14229
rect 1104 14170 22264 14192
rect 1104 14118 4255 14170
rect 4307 14118 4319 14170
rect 4371 14118 4383 14170
rect 4435 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 9545 14170
rect 9597 14118 9609 14170
rect 9661 14118 9673 14170
rect 9725 14118 9737 14170
rect 9789 14118 9801 14170
rect 9853 14118 14835 14170
rect 14887 14118 14899 14170
rect 14951 14118 14963 14170
rect 15015 14118 15027 14170
rect 15079 14118 15091 14170
rect 15143 14118 20125 14170
rect 20177 14118 20189 14170
rect 20241 14118 20253 14170
rect 20305 14118 20317 14170
rect 20369 14118 20381 14170
rect 20433 14118 22264 14170
rect 1104 14096 22264 14118
rect 3970 14056 3976 14068
rect 3344 14028 3976 14056
rect 3142 13880 3148 13932
rect 3200 13880 3206 13932
rect 3344 13929 3372 14028
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 5267 14059 5325 14065
rect 5267 14056 5279 14059
rect 4212 14028 5279 14056
rect 4212 14016 4218 14028
rect 5267 14025 5279 14028
rect 5313 14025 5325 14059
rect 5267 14019 5325 14025
rect 5353 14059 5411 14065
rect 5353 14025 5365 14059
rect 5399 14056 5411 14059
rect 5442 14056 5448 14068
rect 5399 14028 5448 14056
rect 5399 14025 5411 14028
rect 5353 14019 5411 14025
rect 5442 14016 5448 14028
rect 5500 14016 5506 14068
rect 5626 14016 5632 14068
rect 5684 14016 5690 14068
rect 6730 14016 6736 14068
rect 6788 14016 6794 14068
rect 8018 14016 8024 14068
rect 8076 14056 8082 14068
rect 8076 14028 8432 14056
rect 8076 14016 8082 14028
rect 4338 13988 4344 14000
rect 3436 13960 4344 13988
rect 3436 13929 3464 13960
rect 4338 13948 4344 13960
rect 4396 13948 4402 14000
rect 5074 13948 5080 14000
rect 5132 13988 5138 14000
rect 5132 13960 5488 13988
rect 5132 13948 5138 13960
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13889 3479 13923
rect 3677 13923 3735 13929
rect 3677 13920 3689 13923
rect 3421 13883 3479 13889
rect 3528 13892 3689 13920
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13852 3295 13855
rect 3528 13852 3556 13892
rect 3677 13889 3689 13892
rect 3723 13889 3735 13923
rect 3677 13883 3735 13889
rect 5092 13852 5120 13948
rect 5166 13880 5172 13932
rect 5224 13880 5230 13932
rect 5460 13929 5488 13960
rect 5445 13923 5503 13929
rect 5445 13889 5457 13923
rect 5491 13889 5503 13923
rect 5445 13883 5503 13889
rect 5534 13880 5540 13932
rect 5592 13880 5598 13932
rect 5644 13920 5672 14016
rect 6748 13988 6776 14016
rect 8404 13988 8432 14028
rect 8478 14016 8484 14068
rect 8536 14016 8542 14068
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 9953 14059 10011 14065
rect 8720 14028 9352 14056
rect 8720 14016 8726 14028
rect 8573 13991 8631 13997
rect 8573 13988 8585 13991
rect 6564 13960 6776 13988
rect 7116 13960 8340 13988
rect 8404 13960 8585 13988
rect 6564 13929 6592 13960
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 5644 13892 5733 13920
rect 5721 13889 5733 13892
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 6549 13923 6607 13929
rect 6549 13889 6561 13923
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6638 13880 6644 13932
rect 6696 13880 6702 13932
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 7006 13920 7012 13932
rect 6779 13892 7012 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 7006 13880 7012 13892
rect 7064 13880 7070 13932
rect 7116 13929 7144 13960
rect 8312 13932 8340 13960
rect 8573 13957 8585 13960
rect 8619 13957 8631 13991
rect 8573 13951 8631 13957
rect 7374 13929 7380 13932
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 7368 13883 7380 13929
rect 7374 13880 7380 13883
rect 7432 13880 7438 13932
rect 8294 13880 8300 13932
rect 8352 13880 8358 13932
rect 8386 13880 8392 13932
rect 8444 13920 8450 13932
rect 9324 13929 9352 14028
rect 9953 14025 9965 14059
rect 9999 14056 10011 14059
rect 10226 14056 10232 14068
rect 9999 14028 10232 14056
rect 9999 14025 10011 14028
rect 9953 14019 10011 14025
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10870 14016 10876 14068
rect 10928 14016 10934 14068
rect 10962 14016 10968 14068
rect 11020 14056 11026 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 11020 14028 11529 14056
rect 11020 14016 11026 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 12618 14056 12624 14068
rect 11517 14019 11575 14025
rect 12406 14028 12624 14056
rect 9861 13991 9919 13997
rect 9861 13957 9873 13991
rect 9907 13988 9919 13991
rect 10888 13988 10916 14016
rect 11066 13991 11124 13997
rect 11066 13988 11078 13991
rect 9907 13960 10824 13988
rect 10888 13960 11078 13988
rect 9907 13957 9919 13960
rect 9861 13951 9919 13957
rect 10796 13932 10824 13960
rect 11066 13957 11078 13960
rect 11112 13957 11124 13991
rect 12314 13991 12372 13997
rect 11066 13951 11124 13957
rect 11164 13960 11928 13988
rect 8849 13923 8907 13929
rect 8849 13920 8861 13923
rect 8444 13892 8861 13920
rect 8444 13880 8450 13892
rect 8849 13889 8861 13892
rect 8895 13889 8907 13923
rect 8849 13883 8907 13889
rect 9309 13923 9367 13929
rect 9309 13889 9321 13923
rect 9355 13889 9367 13923
rect 10042 13920 10048 13932
rect 9309 13883 9367 13889
rect 9692 13892 10048 13920
rect 3283 13824 3556 13852
rect 4816 13824 5120 13852
rect 5184 13852 5212 13880
rect 5552 13852 5580 13880
rect 5184 13824 5580 13852
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 4816 13793 4844 13824
rect 5810 13812 5816 13864
rect 5868 13812 5874 13864
rect 6822 13852 6828 13864
rect 6104 13824 6828 13852
rect 6104 13793 6132 13824
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 9692 13852 9720 13892
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10778 13880 10784 13932
rect 10836 13920 10842 13932
rect 11164 13920 11192 13960
rect 11900 13929 11928 13960
rect 12314 13957 12326 13991
rect 12360 13988 12372 13991
rect 12406 13988 12434 14028
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 13449 14059 13507 14065
rect 13449 14056 13461 14059
rect 13228 14028 13461 14056
rect 13228 14016 13234 14028
rect 13449 14025 13461 14028
rect 13495 14056 13507 14059
rect 13722 14056 13728 14068
rect 13495 14028 13728 14056
rect 13495 14025 13507 14028
rect 13449 14019 13507 14025
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 14366 14016 14372 14068
rect 14424 14016 14430 14068
rect 14458 14016 14464 14068
rect 14516 14016 14522 14068
rect 15194 14016 15200 14068
rect 15252 14016 15258 14068
rect 15286 14016 15292 14068
rect 15344 14016 15350 14068
rect 15378 14016 15384 14068
rect 15436 14016 15442 14068
rect 15562 14016 15568 14068
rect 15620 14056 15626 14068
rect 16025 14059 16083 14065
rect 16025 14056 16037 14059
rect 15620 14028 16037 14056
rect 15620 14016 15626 14028
rect 16025 14025 16037 14028
rect 16071 14025 16083 14059
rect 16025 14019 16083 14025
rect 16298 14016 16304 14068
rect 16356 14056 16362 14068
rect 16356 14028 16436 14056
rect 16356 14016 16362 14028
rect 12360 13960 12434 13988
rect 12360 13957 12372 13960
rect 12314 13951 12372 13957
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 10836 13892 11192 13920
rect 11624 13892 11713 13920
rect 10836 13880 10842 13892
rect 11624 13864 11652 13892
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 14476 13920 14504 14016
rect 11931 13892 14504 13920
rect 14829 13923 14887 13929
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15212 13920 15240 14016
rect 15304 13988 15332 14016
rect 16408 13997 16436 14028
rect 16942 14016 16948 14068
rect 17000 14016 17006 14068
rect 17497 14059 17555 14065
rect 17497 14025 17509 14059
rect 17543 14056 17555 14059
rect 19058 14056 19064 14068
rect 17543 14028 19064 14056
rect 17543 14025 17555 14028
rect 17497 14019 17555 14025
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 16177 13991 16235 13997
rect 16177 13988 16189 13991
rect 15304 13960 16189 13988
rect 14875 13892 15240 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 15286 13880 15292 13932
rect 15344 13920 15350 13932
rect 15473 13923 15531 13929
rect 15473 13920 15485 13923
rect 15344 13892 15485 13920
rect 15344 13880 15350 13892
rect 15473 13889 15485 13892
rect 15519 13889 15531 13923
rect 15473 13883 15531 13889
rect 15580 13864 15608 13960
rect 16177 13957 16189 13960
rect 16223 13957 16235 13991
rect 16177 13951 16235 13957
rect 16393 13991 16451 13997
rect 16393 13957 16405 13991
rect 16439 13957 16451 13991
rect 16960 13988 16988 14016
rect 16960 13960 17816 13988
rect 16393 13951 16451 13957
rect 8956 13824 9720 13852
rect 8956 13793 8984 13824
rect 11330 13812 11336 13864
rect 11388 13812 11394 13864
rect 11606 13812 11612 13864
rect 11664 13812 11670 13864
rect 12066 13812 12072 13864
rect 12124 13812 12130 13864
rect 14921 13855 14979 13861
rect 14921 13821 14933 13855
rect 14967 13852 14979 13855
rect 15562 13852 15568 13864
rect 14967 13824 15568 13852
rect 14967 13821 14979 13824
rect 14921 13815 14979 13821
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 15933 13855 15991 13861
rect 15933 13821 15945 13855
rect 15979 13852 15991 13855
rect 16408 13852 16436 13951
rect 16758 13880 16764 13932
rect 16816 13920 16822 13932
rect 17788 13929 17816 13960
rect 19996 13960 20576 13988
rect 19996 13932 20024 13960
rect 20548 13932 20576 13960
rect 17313 13923 17371 13929
rect 17313 13920 17325 13923
rect 16816 13892 17325 13920
rect 16816 13880 16822 13892
rect 17313 13889 17325 13892
rect 17359 13889 17371 13923
rect 17313 13883 17371 13889
rect 17773 13923 17831 13929
rect 17773 13889 17785 13923
rect 17819 13889 17831 13923
rect 17773 13883 17831 13889
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13920 18567 13923
rect 18598 13920 18604 13932
rect 18555 13892 18604 13920
rect 18555 13889 18567 13892
rect 18509 13883 18567 13889
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 19978 13880 19984 13932
rect 20036 13880 20042 13932
rect 20254 13929 20260 13932
rect 20248 13920 20260 13929
rect 20215 13892 20260 13920
rect 20248 13883 20260 13892
rect 20254 13880 20260 13883
rect 20312 13880 20318 13932
rect 20530 13880 20536 13932
rect 20588 13880 20594 13932
rect 15979 13824 16436 13852
rect 17129 13855 17187 13861
rect 15979 13821 15991 13824
rect 15933 13815 15991 13821
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17865 13855 17923 13861
rect 17865 13852 17877 13855
rect 17175 13824 17877 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17865 13821 17877 13824
rect 17911 13821 17923 13855
rect 17865 13815 17923 13821
rect 4801 13787 4859 13793
rect 4801 13753 4813 13787
rect 4847 13753 4859 13787
rect 4801 13747 4859 13753
rect 6089 13787 6147 13793
rect 6089 13753 6101 13787
rect 6135 13753 6147 13787
rect 6089 13747 6147 13753
rect 8941 13787 8999 13793
rect 8941 13753 8953 13787
rect 8987 13753 8999 13787
rect 8941 13747 8999 13753
rect 9033 13787 9091 13793
rect 9033 13753 9045 13787
rect 9079 13784 9091 13787
rect 9401 13787 9459 13793
rect 9401 13784 9413 13787
rect 9079 13756 9413 13784
rect 9079 13753 9091 13756
rect 9033 13747 9091 13753
rect 9401 13753 9413 13756
rect 9447 13753 9459 13787
rect 9401 13747 9459 13753
rect 9585 13787 9643 13793
rect 9585 13753 9597 13787
rect 9631 13784 9643 13787
rect 10226 13784 10232 13796
rect 9631 13756 10232 13784
rect 9631 13753 9643 13756
rect 9585 13747 9643 13753
rect 10226 13744 10232 13756
rect 10284 13744 10290 13796
rect 11348 13784 11376 13812
rect 12084 13784 12112 13812
rect 11348 13756 12112 13784
rect 14642 13744 14648 13796
rect 14700 13784 14706 13796
rect 15197 13787 15255 13793
rect 15197 13784 15209 13787
rect 14700 13756 15209 13784
rect 14700 13744 14706 13756
rect 15197 13753 15209 13756
rect 15243 13753 15255 13787
rect 15197 13747 15255 13753
rect 15488 13756 16252 13784
rect 15488 13728 15516 13756
rect 7006 13676 7012 13728
rect 7064 13676 7070 13728
rect 9125 13719 9183 13725
rect 9125 13685 9137 13719
rect 9171 13716 9183 13719
rect 9214 13716 9220 13728
rect 9171 13688 9220 13716
rect 9171 13685 9183 13688
rect 9125 13679 9183 13685
rect 9214 13676 9220 13688
rect 9272 13676 9278 13728
rect 14550 13676 14556 13728
rect 14608 13676 14614 13728
rect 15470 13676 15476 13728
rect 15528 13676 15534 13728
rect 15654 13676 15660 13728
rect 15712 13676 15718 13728
rect 16224 13725 16252 13756
rect 17586 13744 17592 13796
rect 17644 13744 17650 13796
rect 16209 13719 16267 13725
rect 16209 13685 16221 13719
rect 16255 13685 16267 13719
rect 16209 13679 16267 13685
rect 21358 13676 21364 13728
rect 21416 13676 21422 13728
rect 1104 13626 22264 13648
rect 1104 13574 3595 13626
rect 3647 13574 3659 13626
rect 3711 13574 3723 13626
rect 3775 13574 3787 13626
rect 3839 13574 3851 13626
rect 3903 13574 8885 13626
rect 8937 13574 8949 13626
rect 9001 13574 9013 13626
rect 9065 13574 9077 13626
rect 9129 13574 9141 13626
rect 9193 13574 14175 13626
rect 14227 13574 14239 13626
rect 14291 13574 14303 13626
rect 14355 13574 14367 13626
rect 14419 13574 14431 13626
rect 14483 13574 19465 13626
rect 19517 13574 19529 13626
rect 19581 13574 19593 13626
rect 19645 13574 19657 13626
rect 19709 13574 19721 13626
rect 19773 13574 22264 13626
rect 1104 13552 22264 13574
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 8481 13515 8539 13521
rect 8481 13512 8493 13515
rect 7156 13484 8493 13512
rect 7156 13472 7162 13484
rect 8481 13481 8493 13484
rect 8527 13481 8539 13515
rect 8481 13475 8539 13481
rect 9398 13472 9404 13524
rect 9456 13472 9462 13524
rect 10505 13515 10563 13521
rect 10505 13481 10517 13515
rect 10551 13481 10563 13515
rect 10505 13475 10563 13481
rect 15381 13515 15439 13521
rect 15381 13481 15393 13515
rect 15427 13512 15439 13515
rect 15470 13512 15476 13524
rect 15427 13484 15476 13512
rect 15427 13481 15439 13484
rect 15381 13475 15439 13481
rect 9306 13404 9312 13456
rect 9364 13444 9370 13456
rect 9677 13447 9735 13453
rect 9677 13444 9689 13447
rect 9364 13416 9689 13444
rect 9364 13404 9370 13416
rect 9677 13413 9689 13416
rect 9723 13413 9735 13447
rect 10520 13444 10548 13475
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 15562 13472 15568 13524
rect 15620 13472 15626 13524
rect 15654 13472 15660 13524
rect 15712 13472 15718 13524
rect 9677 13407 9735 13413
rect 9784 13416 10548 13444
rect 13541 13447 13599 13453
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 5353 13379 5411 13385
rect 5353 13376 5365 13379
rect 4396 13348 5365 13376
rect 4396 13336 4402 13348
rect 5353 13345 5365 13348
rect 5399 13345 5411 13379
rect 5353 13339 5411 13345
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13376 8999 13379
rect 9214 13376 9220 13388
rect 8987 13348 9220 13376
rect 8987 13345 8999 13348
rect 8941 13339 8999 13345
rect 9214 13336 9220 13348
rect 9272 13376 9278 13388
rect 9784 13376 9812 13416
rect 13541 13413 13553 13447
rect 13587 13413 13599 13447
rect 13541 13407 13599 13413
rect 15197 13447 15255 13453
rect 15197 13413 15209 13447
rect 15243 13444 15255 13447
rect 15580 13444 15608 13472
rect 15243 13416 15608 13444
rect 15243 13413 15255 13416
rect 15197 13407 15255 13413
rect 9272 13348 9812 13376
rect 9272 13336 9278 13348
rect 10226 13336 10232 13388
rect 10284 13336 10290 13388
rect 10502 13336 10508 13388
rect 10560 13376 10566 13388
rect 11057 13379 11115 13385
rect 11057 13376 11069 13379
rect 10560 13348 11069 13376
rect 10560 13336 10566 13348
rect 11057 13345 11069 13348
rect 11103 13345 11115 13379
rect 11057 13339 11115 13345
rect 12066 13336 12072 13388
rect 12124 13376 12130 13388
rect 12161 13379 12219 13385
rect 12161 13376 12173 13379
rect 12124 13348 12173 13376
rect 12124 13336 12130 13348
rect 12161 13345 12173 13348
rect 12207 13345 12219 13379
rect 13556 13376 13584 13407
rect 14553 13379 14611 13385
rect 14553 13376 14565 13379
rect 13556 13348 14565 13376
rect 12161 13339 12219 13345
rect 14553 13345 14565 13348
rect 14599 13345 14611 13379
rect 15672 13376 15700 13472
rect 20533 13379 20591 13385
rect 20533 13376 20545 13379
rect 14553 13339 14611 13345
rect 15304 13348 15700 13376
rect 19536 13348 20545 13376
rect 5620 13311 5678 13317
rect 5620 13277 5632 13311
rect 5666 13308 5678 13311
rect 5994 13308 6000 13320
rect 5666 13280 6000 13308
rect 5666 13277 5678 13280
rect 5620 13271 5678 13277
rect 5994 13268 6000 13280
rect 6052 13268 6058 13320
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 6748 13280 7021 13308
rect 6748 13181 6776 13280
rect 7009 13277 7021 13280
rect 7055 13277 7067 13311
rect 7009 13271 7067 13277
rect 7834 13268 7840 13320
rect 7892 13268 7898 13320
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 8297 13311 8355 13317
rect 8297 13308 8309 13311
rect 8251 13280 8309 13308
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 8297 13277 8309 13280
rect 8343 13277 8355 13311
rect 8297 13271 8355 13277
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13308 10103 13311
rect 10134 13308 10140 13320
rect 10091 13280 10140 13308
rect 10091 13277 10103 13280
rect 10045 13271 10103 13277
rect 10134 13268 10140 13280
rect 10192 13308 10198 13320
rect 15304 13317 15332 13348
rect 10965 13311 11023 13317
rect 10965 13308 10977 13311
rect 10192 13280 10977 13308
rect 10192 13268 10198 13280
rect 10965 13277 10977 13280
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 15289 13311 15347 13317
rect 15289 13277 15301 13311
rect 15335 13277 15347 13311
rect 15473 13311 15531 13317
rect 15473 13308 15485 13311
rect 15289 13271 15347 13277
rect 15396 13280 15485 13308
rect 7466 13200 7472 13252
rect 7524 13240 7530 13252
rect 8021 13243 8079 13249
rect 8021 13240 8033 13243
rect 7524 13212 8033 13240
rect 7524 13200 7530 13212
rect 8021 13209 8033 13212
rect 8067 13209 8079 13243
rect 10778 13240 10784 13252
rect 8021 13203 8079 13209
rect 10152 13212 10784 13240
rect 6733 13175 6791 13181
rect 6733 13141 6745 13175
rect 6779 13141 6791 13175
rect 6733 13135 6791 13141
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 10152 13181 10180 13212
rect 10778 13200 10784 13212
rect 10836 13240 10842 13252
rect 10873 13243 10931 13249
rect 10873 13240 10885 13243
rect 10836 13212 10885 13240
rect 10836 13200 10842 13212
rect 10873 13209 10885 13212
rect 10919 13209 10931 13243
rect 10873 13203 10931 13209
rect 11974 13200 11980 13252
rect 12032 13240 12038 13252
rect 12406 13243 12464 13249
rect 12406 13240 12418 13243
rect 12032 13212 12418 13240
rect 12032 13200 12038 13212
rect 12406 13209 12418 13212
rect 12452 13209 12464 13243
rect 12406 13203 12464 13209
rect 15396 13184 15424 13280
rect 15473 13277 15485 13280
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 17037 13311 17095 13317
rect 17037 13277 17049 13311
rect 17083 13308 17095 13311
rect 17586 13308 17592 13320
rect 17083 13280 17592 13308
rect 17083 13277 17095 13280
rect 17037 13271 17095 13277
rect 17586 13268 17592 13280
rect 17644 13268 17650 13320
rect 18690 13268 18696 13320
rect 18748 13268 18754 13320
rect 19536 13317 19564 13348
rect 20533 13345 20545 13348
rect 20579 13345 20591 13379
rect 20533 13339 20591 13345
rect 18785 13311 18843 13317
rect 18785 13277 18797 13311
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 18969 13311 19027 13317
rect 18969 13277 18981 13311
rect 19015 13308 19027 13311
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 19015 13280 19441 13308
rect 19015 13277 19027 13280
rect 18969 13271 19027 13277
rect 19429 13277 19441 13280
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 19521 13311 19579 13317
rect 19521 13277 19533 13311
rect 19567 13277 19579 13311
rect 19521 13271 19579 13277
rect 20441 13311 20499 13317
rect 20441 13277 20453 13311
rect 20487 13308 20499 13311
rect 20622 13308 20628 13320
rect 20487 13280 20628 13308
rect 20487 13277 20499 13280
rect 20441 13271 20499 13277
rect 16482 13200 16488 13252
rect 16540 13240 16546 13252
rect 16770 13243 16828 13249
rect 16770 13240 16782 13243
rect 16540 13212 16782 13240
rect 16540 13200 16546 13212
rect 16770 13209 16782 13212
rect 16816 13209 16828 13243
rect 16770 13203 16828 13209
rect 18046 13200 18052 13252
rect 18104 13240 18110 13252
rect 18800 13240 18828 13271
rect 20622 13268 20628 13280
rect 20680 13268 20686 13320
rect 20714 13268 20720 13320
rect 20772 13268 20778 13320
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13308 20959 13311
rect 20993 13311 21051 13317
rect 20993 13308 21005 13311
rect 20947 13280 21005 13308
rect 20947 13277 20959 13280
rect 20901 13271 20959 13277
rect 20993 13277 21005 13280
rect 21039 13277 21051 13311
rect 20993 13271 21051 13277
rect 21358 13268 21364 13320
rect 21416 13308 21422 13320
rect 21545 13311 21603 13317
rect 21545 13308 21557 13311
rect 21416 13280 21557 13308
rect 21416 13268 21422 13280
rect 21545 13277 21557 13280
rect 21591 13277 21603 13311
rect 21545 13271 21603 13277
rect 18104 13212 18828 13240
rect 18104 13200 18110 13212
rect 7193 13175 7251 13181
rect 7193 13172 7205 13175
rect 6972 13144 7205 13172
rect 6972 13132 6978 13144
rect 7193 13141 7205 13144
rect 7239 13141 7251 13175
rect 7193 13135 7251 13141
rect 10137 13175 10195 13181
rect 10137 13141 10149 13175
rect 10183 13141 10195 13175
rect 10137 13135 10195 13141
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 14550 13172 14556 13184
rect 13872 13144 14556 13172
rect 13872 13132 13878 13144
rect 14550 13132 14556 13144
rect 14608 13172 14614 13184
rect 14737 13175 14795 13181
rect 14737 13172 14749 13175
rect 14608 13144 14749 13172
rect 14608 13132 14614 13144
rect 14737 13141 14749 13144
rect 14783 13141 14795 13175
rect 14737 13135 14795 13141
rect 14829 13175 14887 13181
rect 14829 13141 14841 13175
rect 14875 13172 14887 13175
rect 15378 13172 15384 13184
rect 14875 13144 15384 13172
rect 14875 13141 14887 13144
rect 14829 13135 14887 13141
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 19242 13132 19248 13184
rect 19300 13132 19306 13184
rect 19702 13132 19708 13184
rect 19760 13132 19766 13184
rect 19794 13132 19800 13184
rect 19852 13132 19858 13184
rect 1104 13082 22264 13104
rect 1104 13030 4255 13082
rect 4307 13030 4319 13082
rect 4371 13030 4383 13082
rect 4435 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 9545 13082
rect 9597 13030 9609 13082
rect 9661 13030 9673 13082
rect 9725 13030 9737 13082
rect 9789 13030 9801 13082
rect 9853 13030 14835 13082
rect 14887 13030 14899 13082
rect 14951 13030 14963 13082
rect 15015 13030 15027 13082
rect 15079 13030 15091 13082
rect 15143 13030 20125 13082
rect 20177 13030 20189 13082
rect 20241 13030 20253 13082
rect 20305 13030 20317 13082
rect 20369 13030 20381 13082
rect 20433 13030 22264 13082
rect 1104 13008 22264 13030
rect 7006 12928 7012 12980
rect 7064 12928 7070 12980
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 7374 12968 7380 12980
rect 7331 12940 7380 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 12989 12971 13047 12977
rect 12989 12968 13001 12971
rect 11848 12940 13001 12968
rect 11848 12928 11854 12940
rect 12989 12937 13001 12940
rect 13035 12968 13047 12971
rect 13035 12940 14688 12968
rect 13035 12937 13047 12940
rect 12989 12931 13047 12937
rect 6822 12860 6828 12912
rect 6880 12860 6886 12912
rect 7024 12900 7052 12928
rect 7024 12872 7420 12900
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 3510 12724 3516 12776
rect 3568 12724 3574 12776
rect 2866 12656 2872 12708
rect 2924 12696 2930 12708
rect 3712 12696 3740 12795
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7009 12835 7067 12841
rect 7009 12832 7021 12835
rect 6972 12804 7021 12832
rect 6972 12792 6978 12804
rect 7009 12801 7021 12804
rect 7055 12801 7067 12835
rect 7009 12795 7067 12801
rect 7098 12792 7104 12844
rect 7156 12792 7162 12844
rect 7392 12841 7420 12872
rect 11698 12860 11704 12912
rect 11756 12860 11762 12912
rect 14550 12860 14556 12912
rect 14608 12860 14614 12912
rect 14660 12900 14688 12940
rect 16482 12928 16488 12980
rect 16540 12928 16546 12980
rect 19705 12971 19763 12977
rect 19705 12937 19717 12971
rect 19751 12968 19763 12971
rect 19978 12968 19984 12980
rect 19751 12940 19984 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 20622 12928 20628 12980
rect 20680 12968 20686 12980
rect 21453 12971 21511 12977
rect 21453 12968 21465 12971
rect 20680 12940 21465 12968
rect 20680 12928 20686 12940
rect 21453 12937 21465 12940
rect 21499 12937 21511 12971
rect 21453 12931 21511 12937
rect 14734 12900 14740 12912
rect 14660 12872 14740 12900
rect 14734 12860 14740 12872
rect 14792 12900 14798 12912
rect 18233 12903 18291 12909
rect 18233 12900 18245 12903
rect 14792 12872 18245 12900
rect 14792 12860 14798 12872
rect 18233 12869 18245 12872
rect 18279 12869 18291 12903
rect 18233 12863 18291 12869
rect 19794 12860 19800 12912
rect 19852 12860 19858 12912
rect 7193 12835 7251 12841
rect 7193 12801 7205 12835
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 14568 12832 14596 12860
rect 15286 12832 15292 12844
rect 14568 12804 15292 12832
rect 7377 12795 7435 12801
rect 4062 12696 4068 12708
rect 2924 12668 4068 12696
rect 2924 12656 2930 12668
rect 4062 12656 4068 12668
rect 4120 12656 4126 12708
rect 6825 12699 6883 12705
rect 6825 12665 6837 12699
rect 6871 12696 6883 12699
rect 7208 12696 7236 12795
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 15654 12792 15660 12844
rect 15712 12792 15718 12844
rect 16022 12792 16028 12844
rect 16080 12792 16086 12844
rect 16209 12835 16267 12841
rect 16209 12801 16221 12835
rect 16255 12832 16267 12835
rect 16301 12835 16359 12841
rect 16301 12832 16313 12835
rect 16255 12804 16313 12832
rect 16255 12801 16267 12804
rect 16209 12795 16267 12801
rect 16301 12801 16313 12804
rect 16347 12801 16359 12835
rect 16301 12795 16359 12801
rect 17957 12835 18015 12841
rect 17957 12801 17969 12835
rect 18003 12832 18015 12835
rect 18046 12832 18052 12844
rect 18003 12804 18052 12832
rect 18003 12801 18015 12804
rect 17957 12795 18015 12801
rect 15378 12724 15384 12776
rect 15436 12724 15442 12776
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12764 15623 12767
rect 15672 12764 15700 12792
rect 15611 12736 15700 12764
rect 15841 12767 15899 12773
rect 15611 12733 15623 12736
rect 15565 12727 15623 12733
rect 15841 12733 15853 12767
rect 15887 12733 15899 12767
rect 16040 12764 16068 12792
rect 17972 12764 18000 12795
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 18141 12835 18199 12841
rect 18141 12801 18153 12835
rect 18187 12832 18199 12835
rect 19812 12832 19840 12860
rect 18187 12804 19840 12832
rect 19996 12832 20024 12928
rect 20073 12835 20131 12841
rect 20073 12832 20085 12835
rect 19996 12804 20085 12832
rect 18187 12801 18199 12804
rect 18141 12795 18199 12801
rect 20073 12801 20085 12804
rect 20119 12801 20131 12835
rect 20329 12835 20387 12841
rect 20329 12832 20341 12835
rect 20073 12795 20131 12801
rect 20180 12804 20341 12832
rect 16040 12736 18000 12764
rect 15841 12727 15899 12733
rect 6871 12668 7236 12696
rect 6871 12665 6883 12668
rect 6825 12659 6883 12665
rect 14642 12656 14648 12708
rect 14700 12696 14706 12708
rect 14921 12699 14979 12705
rect 14921 12696 14933 12699
rect 14700 12668 14933 12696
rect 14700 12656 14706 12668
rect 14921 12665 14933 12668
rect 14967 12665 14979 12699
rect 15396 12696 15424 12724
rect 15856 12696 15884 12727
rect 19702 12724 19708 12776
rect 19760 12764 19766 12776
rect 20180 12764 20208 12804
rect 20329 12801 20341 12804
rect 20375 12801 20387 12835
rect 20329 12795 20387 12801
rect 19760 12736 20208 12764
rect 19760 12724 19766 12736
rect 15396 12668 17908 12696
rect 14921 12659 14979 12665
rect 3881 12631 3939 12637
rect 3881 12597 3893 12631
rect 3927 12628 3939 12631
rect 4430 12628 4436 12640
rect 3927 12600 4436 12628
rect 3927 12597 3939 12600
rect 3881 12591 3939 12597
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 17494 12588 17500 12640
rect 17552 12628 17558 12640
rect 17773 12631 17831 12637
rect 17773 12628 17785 12631
rect 17552 12600 17785 12628
rect 17552 12588 17558 12600
rect 17773 12597 17785 12600
rect 17819 12597 17831 12631
rect 17880 12628 17908 12668
rect 21450 12628 21456 12640
rect 17880 12600 21456 12628
rect 17773 12591 17831 12597
rect 21450 12588 21456 12600
rect 21508 12588 21514 12640
rect 1104 12538 22264 12560
rect 1104 12486 3595 12538
rect 3647 12486 3659 12538
rect 3711 12486 3723 12538
rect 3775 12486 3787 12538
rect 3839 12486 3851 12538
rect 3903 12486 8885 12538
rect 8937 12486 8949 12538
rect 9001 12486 9013 12538
rect 9065 12486 9077 12538
rect 9129 12486 9141 12538
rect 9193 12486 14175 12538
rect 14227 12486 14239 12538
rect 14291 12486 14303 12538
rect 14355 12486 14367 12538
rect 14419 12486 14431 12538
rect 14483 12486 19465 12538
rect 19517 12486 19529 12538
rect 19581 12486 19593 12538
rect 19645 12486 19657 12538
rect 19709 12486 19721 12538
rect 19773 12486 22264 12538
rect 1104 12464 22264 12486
rect 3510 12384 3516 12436
rect 3568 12424 3574 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3568 12396 3801 12424
rect 3568 12384 3574 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3789 12387 3847 12393
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 5810 12424 5816 12436
rect 5592 12396 5816 12424
rect 5592 12384 5598 12396
rect 5810 12384 5816 12396
rect 5868 12424 5874 12436
rect 10410 12424 10416 12436
rect 5868 12396 10416 12424
rect 5868 12384 5874 12396
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 10502 12384 10508 12436
rect 10560 12384 10566 12436
rect 11974 12384 11980 12436
rect 12032 12384 12038 12436
rect 17586 12384 17592 12436
rect 17644 12424 17650 12436
rect 19978 12424 19984 12436
rect 17644 12396 19984 12424
rect 17644 12384 17650 12396
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20714 12424 20720 12436
rect 20180 12396 20720 12424
rect 3418 12316 3424 12368
rect 3476 12356 3482 12368
rect 3476 12328 3740 12356
rect 3476 12316 3482 12328
rect 3712 12288 3740 12328
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 4120 12328 5764 12356
rect 4120 12316 4126 12328
rect 4341 12291 4399 12297
rect 4341 12288 4353 12291
rect 3712 12260 4353 12288
rect 4341 12257 4353 12260
rect 4387 12257 4399 12291
rect 4341 12251 4399 12257
rect 5736 12232 5764 12328
rect 13814 12288 13820 12300
rect 10888 12260 13820 12288
rect 1578 12180 1584 12232
rect 1636 12220 1642 12232
rect 2041 12223 2099 12229
rect 2041 12220 2053 12223
rect 1636 12192 2053 12220
rect 1636 12180 1642 12192
rect 2041 12189 2053 12192
rect 2087 12220 2099 12223
rect 4154 12220 4160 12232
rect 2087 12192 4160 12220
rect 2087 12189 2099 12192
rect 2041 12183 2099 12189
rect 4154 12180 4160 12192
rect 4212 12180 4218 12232
rect 4430 12180 4436 12232
rect 4488 12220 4494 12232
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 4488 12192 4721 12220
rect 4488 12180 4494 12192
rect 4709 12189 4721 12192
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 5258 12180 5264 12232
rect 5316 12180 5322 12232
rect 5534 12180 5540 12232
rect 5592 12180 5598 12232
rect 5718 12180 5724 12232
rect 5776 12180 5782 12232
rect 5905 12223 5963 12229
rect 5905 12189 5917 12223
rect 5951 12220 5963 12223
rect 6181 12223 6239 12229
rect 6181 12220 6193 12223
rect 5951 12192 6193 12220
rect 5951 12189 5963 12192
rect 5905 12183 5963 12189
rect 6181 12189 6193 12192
rect 6227 12189 6239 12223
rect 6181 12183 6239 12189
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12220 9183 12223
rect 9950 12220 9956 12232
rect 9171 12192 9956 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 10888 12229 10916 12260
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 17604 12297 17632 12384
rect 18690 12316 18696 12368
rect 18748 12356 18754 12368
rect 19245 12359 19303 12365
rect 19245 12356 19257 12359
rect 18748 12328 19257 12356
rect 18748 12316 18754 12328
rect 19245 12325 19257 12328
rect 19291 12325 19303 12359
rect 19245 12319 19303 12325
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12257 17647 12291
rect 17589 12251 17647 12257
rect 10873 12223 10931 12229
rect 10873 12220 10885 12223
rect 10704 12192 10885 12220
rect 2130 12112 2136 12164
rect 2188 12152 2194 12164
rect 2286 12155 2344 12161
rect 2286 12152 2298 12155
rect 2188 12124 2298 12152
rect 2188 12112 2194 12124
rect 2286 12121 2298 12124
rect 2332 12121 2344 12155
rect 2286 12115 2344 12121
rect 9392 12155 9450 12161
rect 9392 12121 9404 12155
rect 9438 12152 9450 12155
rect 10318 12152 10324 12164
rect 9438 12124 10324 12152
rect 9438 12121 9450 12124
rect 9392 12115 9450 12121
rect 10318 12112 10324 12124
rect 10376 12112 10382 12164
rect 4525 12087 4583 12093
rect 4525 12053 4537 12087
rect 4571 12084 4583 12087
rect 4614 12084 4620 12096
rect 4571 12056 4620 12084
rect 4571 12053 4583 12056
rect 4525 12047 4583 12053
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 4890 12044 4896 12096
rect 4948 12084 4954 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 4948 12056 5089 12084
rect 4948 12044 4954 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5077 12047 5135 12053
rect 5994 12044 6000 12096
rect 6052 12044 6058 12096
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 10704 12084 10732 12192
rect 10873 12189 10885 12192
rect 10919 12189 10931 12223
rect 10873 12183 10931 12189
rect 11057 12223 11115 12229
rect 11057 12189 11069 12223
rect 11103 12189 11115 12223
rect 11057 12183 11115 12189
rect 11241 12223 11299 12229
rect 11241 12189 11253 12223
rect 11287 12220 11299 12223
rect 11793 12223 11851 12229
rect 11793 12220 11805 12223
rect 11287 12192 11805 12220
rect 11287 12189 11299 12192
rect 11241 12183 11299 12189
rect 11793 12189 11805 12192
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12220 14519 12223
rect 14550 12220 14556 12232
rect 14507 12192 14556 12220
rect 14507 12189 14519 12192
rect 14461 12183 14519 12189
rect 11072 12152 11100 12183
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 17310 12180 17316 12232
rect 17368 12180 17374 12232
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 18984 12192 19809 12220
rect 15930 12152 15936 12164
rect 10796 12124 11100 12152
rect 12406 12124 15936 12152
rect 10796 12096 10824 12124
rect 8720 12056 10732 12084
rect 8720 12044 8726 12056
rect 10778 12044 10784 12096
rect 10836 12044 10842 12096
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 11882 12084 11888 12096
rect 11296 12056 11888 12084
rect 11296 12044 11302 12056
rect 11882 12044 11888 12056
rect 11940 12084 11946 12096
rect 12406 12084 12434 12124
rect 15930 12112 15936 12124
rect 15988 12112 15994 12164
rect 17834 12155 17892 12161
rect 17834 12152 17846 12155
rect 17512 12124 17846 12152
rect 11940 12056 12434 12084
rect 11940 12044 11946 12056
rect 12986 12044 12992 12096
rect 13044 12084 13050 12096
rect 13906 12084 13912 12096
rect 13044 12056 13912 12084
rect 13044 12044 13050 12056
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 17512 12093 17540 12124
rect 17834 12121 17846 12124
rect 17880 12121 17892 12155
rect 17834 12115 17892 12121
rect 18984 12093 19012 12192
rect 19797 12189 19809 12192
rect 19843 12220 19855 12223
rect 19886 12220 19892 12232
rect 19843 12192 19892 12220
rect 19843 12189 19855 12192
rect 19797 12183 19855 12189
rect 19886 12180 19892 12192
rect 19944 12180 19950 12232
rect 20180 12229 20208 12396
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 21450 12384 21456 12436
rect 21508 12384 21514 12436
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12189 20223 12223
rect 20165 12183 20223 12189
rect 20349 12223 20407 12229
rect 20349 12189 20361 12223
rect 20395 12189 20407 12223
rect 20349 12183 20407 12189
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12189 20499 12223
rect 20441 12183 20499 12189
rect 14277 12087 14335 12093
rect 14277 12084 14289 12087
rect 14056 12056 14289 12084
rect 14056 12044 14062 12056
rect 14277 12053 14289 12056
rect 14323 12053 14335 12087
rect 14277 12047 14335 12053
rect 17497 12087 17555 12093
rect 17497 12053 17509 12087
rect 17543 12053 17555 12087
rect 17497 12047 17555 12053
rect 18969 12087 19027 12093
rect 18969 12053 18981 12087
rect 19015 12053 19027 12087
rect 18969 12047 19027 12053
rect 19150 12044 19156 12096
rect 19208 12084 19214 12096
rect 19981 12087 20039 12093
rect 19981 12084 19993 12087
rect 19208 12056 19993 12084
rect 19208 12044 19214 12056
rect 19981 12053 19993 12056
rect 20027 12053 20039 12087
rect 20364 12084 20392 12183
rect 20456 12152 20484 12183
rect 20714 12180 20720 12232
rect 20772 12180 20778 12232
rect 20990 12152 20996 12164
rect 20456 12124 20996 12152
rect 20990 12112 20996 12124
rect 21048 12112 21054 12164
rect 20530 12084 20536 12096
rect 20364 12056 20536 12084
rect 19981 12047 20039 12053
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 1104 11994 22264 12016
rect 1104 11942 4255 11994
rect 4307 11942 4319 11994
rect 4371 11942 4383 11994
rect 4435 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 9545 11994
rect 9597 11942 9609 11994
rect 9661 11942 9673 11994
rect 9725 11942 9737 11994
rect 9789 11942 9801 11994
rect 9853 11942 14835 11994
rect 14887 11942 14899 11994
rect 14951 11942 14963 11994
rect 15015 11942 15027 11994
rect 15079 11942 15091 11994
rect 15143 11942 20125 11994
rect 20177 11942 20189 11994
rect 20241 11942 20253 11994
rect 20305 11942 20317 11994
rect 20369 11942 20381 11994
rect 20433 11942 22264 11994
rect 1104 11920 22264 11942
rect 4614 11840 4620 11892
rect 4672 11840 4678 11892
rect 5534 11840 5540 11892
rect 5592 11840 5598 11892
rect 8662 11840 8668 11892
rect 8720 11840 8726 11892
rect 9674 11880 9680 11892
rect 9416 11852 9680 11880
rect 4332 11815 4390 11821
rect 4332 11781 4344 11815
rect 4378 11812 4390 11815
rect 4632 11812 4660 11840
rect 4378 11784 4660 11812
rect 4378 11781 4390 11784
rect 4332 11775 4390 11781
rect 6362 11772 6368 11824
rect 6420 11772 6426 11824
rect 6581 11815 6639 11821
rect 6581 11781 6593 11815
rect 6627 11812 6639 11815
rect 6730 11812 6736 11824
rect 6627 11784 6736 11812
rect 6627 11781 6639 11784
rect 6581 11775 6639 11781
rect 6730 11772 6736 11784
rect 6788 11772 6794 11824
rect 9416 11821 9444 11852
rect 9674 11840 9680 11852
rect 9732 11880 9738 11892
rect 10226 11880 10232 11892
rect 9732 11852 10232 11880
rect 9732 11840 9738 11852
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 10318 11840 10324 11892
rect 10376 11840 10382 11892
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 12986 11880 12992 11892
rect 10928 11852 12992 11880
rect 10928 11840 10934 11852
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 15565 11883 15623 11889
rect 13096 11852 14228 11880
rect 9401 11815 9459 11821
rect 9401 11781 9413 11815
rect 9447 11781 9459 11815
rect 10134 11812 10140 11824
rect 9401 11775 9459 11781
rect 9968 11784 10140 11812
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11744 1547 11747
rect 1578 11744 1584 11756
rect 1535 11716 1584 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 1762 11753 1768 11756
rect 1756 11707 1768 11753
rect 1762 11704 1768 11707
rect 1820 11704 1826 11756
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11744 4123 11747
rect 4154 11744 4160 11756
rect 4111 11716 4160 11744
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 4154 11704 4160 11716
rect 4212 11704 4218 11756
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11713 6975 11747
rect 6917 11707 6975 11713
rect 3697 11679 3755 11685
rect 3697 11645 3709 11679
rect 3743 11645 3755 11679
rect 3697 11639 3755 11645
rect 2869 11611 2927 11617
rect 2869 11577 2881 11611
rect 2915 11608 2927 11611
rect 3326 11608 3332 11620
rect 2915 11580 3332 11608
rect 2915 11577 2927 11580
rect 2869 11571 2927 11577
rect 3326 11568 3332 11580
rect 3384 11608 3390 11620
rect 3712 11608 3740 11639
rect 6178 11636 6184 11688
rect 6236 11636 6242 11688
rect 6932 11608 6960 11707
rect 7098 11704 7104 11756
rect 7156 11704 7162 11756
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11744 7435 11747
rect 7929 11747 7987 11753
rect 7929 11744 7941 11747
rect 7423 11716 7941 11744
rect 7423 11713 7435 11716
rect 7377 11707 7435 11713
rect 7929 11713 7941 11716
rect 7975 11744 7987 11747
rect 8018 11744 8024 11756
rect 7975 11716 8024 11744
rect 7975 11713 7987 11716
rect 7929 11707 7987 11713
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 9968 11753 9996 11784
rect 10134 11772 10140 11784
rect 10192 11812 10198 11824
rect 10192 11784 13032 11812
rect 10192 11772 10198 11784
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10045 11747 10103 11753
rect 10045 11713 10057 11747
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11744 10287 11747
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 10275 11716 10517 11744
rect 10275 11713 10287 11716
rect 10229 11707 10287 11713
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11676 7619 11679
rect 7653 11679 7711 11685
rect 7653 11676 7665 11679
rect 7607 11648 7665 11676
rect 7607 11645 7619 11648
rect 7561 11639 7619 11645
rect 7653 11645 7665 11648
rect 7699 11645 7711 11679
rect 7653 11639 7711 11645
rect 9766 11636 9772 11688
rect 9824 11676 9830 11688
rect 10060 11676 10088 11707
rect 10778 11704 10784 11756
rect 10836 11704 10842 11756
rect 11330 11704 11336 11756
rect 11388 11704 11394 11756
rect 12526 11704 12532 11756
rect 12584 11704 12590 11756
rect 12894 11704 12900 11756
rect 12952 11704 12958 11756
rect 10796 11676 10824 11704
rect 9824 11648 10824 11676
rect 10965 11679 11023 11685
rect 9824 11636 9830 11648
rect 10965 11645 10977 11679
rect 11011 11645 11023 11679
rect 10965 11639 11023 11645
rect 3384 11580 3740 11608
rect 5000 11580 6960 11608
rect 9677 11611 9735 11617
rect 3384 11568 3390 11580
rect 3050 11500 3056 11552
rect 3108 11540 3114 11552
rect 3145 11543 3203 11549
rect 3145 11540 3157 11543
rect 3108 11512 3157 11540
rect 3108 11500 3114 11512
rect 3145 11509 3157 11512
rect 3191 11509 3203 11543
rect 3145 11503 3203 11509
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 5000 11540 5028 11580
rect 9677 11577 9689 11611
rect 9723 11608 9735 11611
rect 10410 11608 10416 11620
rect 9723 11580 10416 11608
rect 9723 11577 9735 11580
rect 9677 11571 9735 11577
rect 10410 11568 10416 11580
rect 10468 11568 10474 11620
rect 10980 11608 11008 11639
rect 12250 11636 12256 11688
rect 12308 11636 12314 11688
rect 12802 11608 12808 11620
rect 10980 11580 12808 11608
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 4304 11512 5028 11540
rect 5445 11543 5503 11549
rect 4304 11500 4310 11512
rect 5445 11509 5457 11543
rect 5491 11540 5503 11543
rect 5902 11540 5908 11552
rect 5491 11512 5908 11540
rect 5491 11509 5503 11512
rect 5445 11503 5503 11509
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6546 11500 6552 11552
rect 6604 11500 6610 11552
rect 6733 11543 6791 11549
rect 6733 11509 6745 11543
rect 6779 11540 6791 11543
rect 7282 11540 7288 11552
rect 6779 11512 7288 11540
rect 6779 11509 6791 11512
rect 6733 11503 6791 11509
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 10594 11500 10600 11552
rect 10652 11500 10658 11552
rect 11146 11500 11152 11552
rect 11204 11500 11210 11552
rect 11609 11543 11667 11549
rect 11609 11509 11621 11543
rect 11655 11540 11667 11543
rect 11790 11540 11796 11552
rect 11655 11512 11796 11540
rect 11655 11509 11667 11512
rect 11609 11503 11667 11509
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 12342 11500 12348 11552
rect 12400 11500 12406 11552
rect 13004 11540 13032 11784
rect 13096 11753 13124 11852
rect 13998 11812 14004 11824
rect 13924 11784 14004 11812
rect 13924 11753 13952 11784
rect 13998 11772 14004 11784
rect 14056 11772 14062 11824
rect 14200 11812 14228 11852
rect 15565 11849 15577 11883
rect 15611 11880 15623 11883
rect 15746 11880 15752 11892
rect 15611 11852 15752 11880
rect 15611 11849 15623 11852
rect 15565 11843 15623 11849
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 20165 11883 20223 11889
rect 15856 11852 19380 11880
rect 14642 11812 14648 11824
rect 14200 11784 14648 11812
rect 14642 11772 14648 11784
rect 14700 11772 14706 11824
rect 15856 11753 15884 11852
rect 15930 11772 15936 11824
rect 15988 11772 15994 11824
rect 16758 11772 16764 11824
rect 16816 11772 16822 11824
rect 18316 11815 18374 11821
rect 18316 11781 18328 11815
rect 18362 11812 18374 11815
rect 19242 11812 19248 11824
rect 18362 11784 19248 11812
rect 18362 11781 18374 11784
rect 18316 11775 18374 11781
rect 19242 11772 19248 11784
rect 19300 11772 19306 11824
rect 19352 11812 19380 11852
rect 20165 11849 20177 11883
rect 20211 11880 20223 11883
rect 20530 11880 20536 11892
rect 20211 11852 20536 11880
rect 20211 11849 20223 11852
rect 20165 11843 20223 11849
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 20714 11840 20720 11892
rect 20772 11880 20778 11892
rect 21085 11883 21143 11889
rect 21085 11880 21097 11883
rect 20772 11852 21097 11880
rect 20772 11840 20778 11852
rect 21085 11849 21097 11852
rect 21131 11849 21143 11883
rect 21085 11843 21143 11849
rect 19352 11784 20484 11812
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11744 13415 11747
rect 13909 11747 13967 11753
rect 13909 11744 13921 11747
rect 13403 11716 13921 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13909 11713 13921 11716
rect 13955 11713 13967 11747
rect 13909 11707 13967 11713
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11744 15255 11747
rect 15657 11747 15715 11753
rect 15657 11744 15669 11747
rect 15243 11716 15669 11744
rect 15243 11713 15255 11716
rect 15197 11707 15255 11713
rect 15657 11713 15669 11716
rect 15703 11744 15715 11747
rect 15841 11747 15899 11753
rect 15841 11744 15853 11747
rect 15703 11716 15853 11744
rect 15703 11713 15715 11716
rect 15657 11707 15715 11713
rect 15841 11713 15853 11716
rect 15887 11713 15899 11747
rect 15841 11707 15899 11713
rect 16022 11704 16028 11756
rect 16080 11744 16086 11756
rect 16301 11747 16359 11753
rect 16301 11744 16313 11747
rect 16080 11716 16313 11744
rect 16080 11704 16086 11716
rect 16301 11713 16313 11716
rect 16347 11744 16359 11747
rect 16776 11744 16804 11772
rect 16347 11716 16804 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 17586 11704 17592 11756
rect 17644 11744 17650 11756
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 17644 11716 18061 11744
rect 17644 11704 17650 11716
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 18049 11707 18107 11713
rect 19444 11716 20361 11744
rect 13541 11679 13599 11685
rect 13541 11645 13553 11679
rect 13587 11676 13599 11679
rect 13633 11679 13691 11685
rect 13633 11676 13645 11679
rect 13587 11648 13645 11676
rect 13587 11645 13599 11648
rect 13541 11639 13599 11645
rect 13633 11645 13645 11648
rect 13679 11645 13691 11679
rect 13633 11639 13691 11645
rect 14366 11636 14372 11688
rect 14424 11676 14430 11688
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 14424 11648 14933 11676
rect 14424 11636 14430 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11676 16175 11679
rect 16669 11679 16727 11685
rect 16669 11676 16681 11679
rect 16163 11648 16681 11676
rect 16163 11645 16175 11648
rect 16117 11639 16175 11645
rect 16669 11645 16681 11648
rect 16715 11645 16727 11679
rect 16669 11639 16727 11645
rect 17218 11636 17224 11688
rect 17276 11636 17282 11688
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 19444 11676 19472 11716
rect 20349 11713 20361 11716
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 19300 11648 19472 11676
rect 19613 11679 19671 11685
rect 19300 11636 19306 11648
rect 19613 11645 19625 11679
rect 19659 11676 19671 11679
rect 19659 11648 19840 11676
rect 19659 11645 19671 11648
rect 19613 11639 19671 11645
rect 14645 11611 14703 11617
rect 14645 11577 14657 11611
rect 14691 11577 14703 11611
rect 14645 11571 14703 11577
rect 14660 11540 14688 11571
rect 19812 11552 19840 11648
rect 20456 11608 20484 11784
rect 20533 11747 20591 11753
rect 20533 11713 20545 11747
rect 20579 11713 20591 11747
rect 20732 11744 20760 11840
rect 20990 11772 20996 11824
rect 21048 11772 21054 11824
rect 20809 11747 20867 11753
rect 20809 11744 20821 11747
rect 20732 11716 20821 11744
rect 20533 11707 20591 11713
rect 20809 11713 20821 11716
rect 20855 11713 20867 11747
rect 20809 11707 20867 11713
rect 20548 11676 20576 11707
rect 21266 11704 21272 11756
rect 21324 11704 21330 11756
rect 21637 11747 21695 11753
rect 21637 11713 21649 11747
rect 21683 11713 21695 11747
rect 21637 11707 21695 11713
rect 20714 11676 20720 11688
rect 20548 11648 20720 11676
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 21652 11676 21680 11707
rect 22186 11676 22192 11688
rect 21652 11648 22192 11676
rect 22186 11636 22192 11648
rect 22244 11636 22250 11688
rect 21453 11611 21511 11617
rect 21453 11608 21465 11611
rect 20456 11580 21465 11608
rect 21453 11577 21465 11580
rect 21499 11577 21511 11611
rect 21453 11571 21511 11577
rect 13004 11512 14688 11540
rect 16482 11500 16488 11552
rect 16540 11500 16546 11552
rect 19429 11543 19487 11549
rect 19429 11509 19441 11543
rect 19475 11540 19487 11543
rect 19794 11540 19800 11552
rect 19475 11512 19800 11540
rect 19475 11509 19487 11512
rect 19429 11503 19487 11509
rect 19794 11500 19800 11512
rect 19852 11500 19858 11552
rect 1104 11450 22264 11472
rect 1104 11398 3595 11450
rect 3647 11398 3659 11450
rect 3711 11398 3723 11450
rect 3775 11398 3787 11450
rect 3839 11398 3851 11450
rect 3903 11398 8885 11450
rect 8937 11398 8949 11450
rect 9001 11398 9013 11450
rect 9065 11398 9077 11450
rect 9129 11398 9141 11450
rect 9193 11398 14175 11450
rect 14227 11398 14239 11450
rect 14291 11398 14303 11450
rect 14355 11398 14367 11450
rect 14419 11398 14431 11450
rect 14483 11398 19465 11450
rect 19517 11398 19529 11450
rect 19581 11398 19593 11450
rect 19645 11398 19657 11450
rect 19709 11398 19721 11450
rect 19773 11398 22264 11450
rect 1104 11376 22264 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1762 11336 1768 11348
rect 1719 11308 1768 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 2130 11296 2136 11348
rect 2188 11296 2194 11348
rect 2866 11336 2872 11348
rect 2746 11308 2872 11336
rect 2225 11203 2283 11209
rect 2225 11200 2237 11203
rect 1872 11172 2237 11200
rect 1872 11141 1900 11172
rect 2225 11169 2237 11172
rect 2271 11169 2283 11203
rect 2746 11200 2774 11308
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3050 11296 3056 11348
rect 3108 11296 3114 11348
rect 3418 11296 3424 11348
rect 3476 11296 3482 11348
rect 4246 11336 4252 11348
rect 3620 11308 4252 11336
rect 3068 11209 3096 11296
rect 3620 11277 3648 11308
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 4341 11339 4399 11345
rect 4341 11305 4353 11339
rect 4387 11336 4399 11339
rect 6546 11336 6552 11348
rect 4387 11308 6552 11336
rect 4387 11305 4399 11308
rect 4341 11299 4399 11305
rect 6546 11296 6552 11308
rect 6604 11296 6610 11348
rect 9766 11336 9772 11348
rect 7484 11308 9772 11336
rect 3605 11271 3663 11277
rect 3605 11237 3617 11271
rect 3651 11237 3663 11271
rect 3605 11231 3663 11237
rect 6362 11228 6368 11280
rect 6420 11268 6426 11280
rect 6638 11268 6644 11280
rect 6420 11240 6644 11268
rect 6420 11228 6426 11240
rect 6638 11228 6644 11240
rect 6696 11268 6702 11280
rect 7101 11271 7159 11277
rect 7101 11268 7113 11271
rect 6696 11240 7113 11268
rect 6696 11228 6702 11240
rect 7101 11237 7113 11240
rect 7147 11237 7159 11271
rect 7101 11231 7159 11237
rect 3053 11203 3111 11209
rect 2225 11163 2283 11169
rect 2424 11172 3004 11200
rect 2424 11144 2452 11172
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11101 1915 11135
rect 1857 11095 1915 11101
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11101 2007 11135
rect 1949 11095 2007 11101
rect 1964 11064 1992 11095
rect 2406 11092 2412 11144
rect 2464 11092 2470 11144
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11132 2651 11135
rect 2774 11132 2780 11144
rect 2639 11104 2780 11132
rect 2639 11101 2651 11104
rect 2593 11095 2651 11101
rect 2774 11092 2780 11104
rect 2832 11092 2838 11144
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 2976 11132 3004 11172
rect 3053 11169 3065 11203
rect 3099 11169 3111 11203
rect 3053 11163 3111 11169
rect 3344 11172 4108 11200
rect 3344 11141 3372 11172
rect 3329 11135 3387 11141
rect 3329 11132 3341 11135
rect 2915 11104 3004 11132
rect 3068 11104 3341 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 2685 11067 2743 11073
rect 2685 11064 2697 11067
rect 1964 11036 2697 11064
rect 2685 11033 2697 11036
rect 2731 11033 2743 11067
rect 2685 11027 2743 11033
rect 2958 10956 2964 11008
rect 3016 10996 3022 11008
rect 3068 10996 3096 11104
rect 3329 11101 3341 11104
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 3418 11092 3424 11144
rect 3476 11092 3482 11144
rect 3510 11092 3516 11144
rect 3568 11132 3574 11144
rect 4080 11141 4108 11172
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4614 11200 4620 11212
rect 4212 11172 4620 11200
rect 4212 11160 4218 11172
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 7484 11200 7512 11308
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 10594 11336 10600 11348
rect 10336 11308 10600 11336
rect 8754 11228 8760 11280
rect 8812 11268 8818 11280
rect 9217 11271 9275 11277
rect 9217 11268 9229 11271
rect 8812 11240 9229 11268
rect 8812 11228 8818 11240
rect 9217 11237 9229 11240
rect 9263 11237 9275 11271
rect 9217 11231 9275 11237
rect 6880 11172 7512 11200
rect 6880 11160 6886 11172
rect 4890 11141 4896 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3568 11104 3985 11132
rect 3568 11092 3574 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 4884 11132 4896 11141
rect 4851 11104 4896 11132
rect 4065 11095 4123 11101
rect 4884 11095 4896 11104
rect 4890 11092 4896 11095
rect 4948 11092 4954 11144
rect 6362 11092 6368 11144
rect 6420 11092 6426 11144
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11132 8539 11135
rect 9950 11132 9956 11144
rect 8527 11104 9956 11132
rect 8527 11101 8539 11104
rect 8481 11095 8539 11101
rect 9950 11092 9956 11104
rect 10008 11092 10014 11144
rect 10336 11141 10364 11308
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 11793 11339 11851 11345
rect 11793 11305 11805 11339
rect 11839 11336 11851 11339
rect 12618 11336 12624 11348
rect 11839 11308 12624 11336
rect 11839 11305 11851 11308
rect 11793 11299 11851 11305
rect 12618 11296 12624 11308
rect 12676 11336 12682 11348
rect 13909 11339 13967 11345
rect 12676 11308 13400 11336
rect 12676 11296 12682 11308
rect 13372 11277 13400 11308
rect 13909 11305 13921 11339
rect 13955 11336 13967 11339
rect 14461 11339 14519 11345
rect 14461 11336 14473 11339
rect 13955 11308 14473 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 14461 11305 14473 11308
rect 14507 11305 14519 11339
rect 14461 11299 14519 11305
rect 14550 11296 14556 11348
rect 14608 11296 14614 11348
rect 14642 11296 14648 11348
rect 14700 11336 14706 11348
rect 14737 11339 14795 11345
rect 14737 11336 14749 11339
rect 14700 11308 14749 11336
rect 14700 11296 14706 11308
rect 14737 11305 14749 11308
rect 14783 11305 14795 11339
rect 15197 11339 15255 11345
rect 15197 11336 15209 11339
rect 14737 11299 14795 11305
rect 14844 11308 15209 11336
rect 13265 11271 13323 11277
rect 13265 11237 13277 11271
rect 13311 11237 13323 11271
rect 13265 11231 13323 11237
rect 13357 11271 13415 11277
rect 13357 11237 13369 11271
rect 13403 11237 13415 11271
rect 13357 11231 13415 11237
rect 14277 11271 14335 11277
rect 14277 11237 14289 11271
rect 14323 11268 14335 11271
rect 14568 11268 14596 11296
rect 14323 11240 14596 11268
rect 14323 11237 14335 11240
rect 14277 11231 14335 11237
rect 13280 11200 13308 11231
rect 13538 11200 13544 11212
rect 13280 11172 13544 11200
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11132 10471 11135
rect 10962 11132 10968 11144
rect 10459 11104 10968 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 10962 11092 10968 11104
rect 11020 11132 11026 11144
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 11020 11104 11897 11132
rect 11020 11092 11026 11104
rect 11885 11101 11897 11104
rect 11931 11132 11943 11135
rect 11931 11104 13860 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 3145 11067 3203 11073
rect 3145 11033 3157 11067
rect 3191 11033 3203 11067
rect 3145 11027 3203 11033
rect 3016 10968 3096 10996
rect 3160 10996 3188 11027
rect 3326 10996 3332 11008
rect 3160 10968 3332 10996
rect 3016 10956 3022 10968
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 3436 10996 3464 11092
rect 3789 11067 3847 11073
rect 3789 11033 3801 11067
rect 3835 11033 3847 11067
rect 4157 11067 4215 11073
rect 4157 11064 4169 11067
rect 3789 11027 3847 11033
rect 3896 11036 4169 11064
rect 3804 10996 3832 11027
rect 3896 11008 3924 11036
rect 4157 11033 4169 11036
rect 4203 11033 4215 11067
rect 4157 11027 4215 11033
rect 7742 11024 7748 11076
rect 7800 11064 7806 11076
rect 8214 11067 8272 11073
rect 8214 11064 8226 11067
rect 7800 11036 8226 11064
rect 7800 11024 7806 11036
rect 8214 11033 8226 11036
rect 8260 11033 8272 11067
rect 8214 11027 8272 11033
rect 9033 11067 9091 11073
rect 9033 11033 9045 11067
rect 9079 11064 9091 11067
rect 9582 11064 9588 11076
rect 9079 11036 9588 11064
rect 9079 11033 9091 11036
rect 9033 11027 9091 11033
rect 9582 11024 9588 11036
rect 9640 11024 9646 11076
rect 9677 11067 9735 11073
rect 9677 11033 9689 11067
rect 9723 11064 9735 11067
rect 10680 11067 10738 11073
rect 9723 11036 10640 11064
rect 9723 11033 9735 11036
rect 9677 11027 9735 11033
rect 3436 10968 3832 10996
rect 3878 10956 3884 11008
rect 3936 10956 3942 11008
rect 5997 10999 6055 11005
rect 5997 10965 6009 10999
rect 6043 10996 6055 10999
rect 6178 10996 6184 11008
rect 6043 10968 6184 10996
rect 6043 10965 6055 10968
rect 5997 10959 6055 10965
rect 6178 10956 6184 10968
rect 6236 10996 6242 11008
rect 6546 10996 6552 11008
rect 6236 10968 6552 10996
rect 6236 10956 6242 10968
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 7006 10956 7012 11008
rect 7064 10956 7070 11008
rect 10134 10956 10140 11008
rect 10192 10956 10198 11008
rect 10612 10996 10640 11036
rect 10680 11033 10692 11067
rect 10726 11064 10738 11067
rect 11146 11064 11152 11076
rect 10726 11036 11152 11064
rect 10726 11033 10738 11036
rect 10680 11027 10738 11033
rect 11146 11024 11152 11036
rect 11204 11024 11210 11076
rect 11238 11024 11244 11076
rect 11296 11024 11302 11076
rect 12152 11067 12210 11073
rect 12152 11033 12164 11067
rect 12198 11064 12210 11067
rect 12342 11064 12348 11076
rect 12198 11036 12348 11064
rect 12198 11033 12210 11036
rect 12152 11027 12210 11033
rect 12342 11024 12348 11036
rect 12400 11024 12406 11076
rect 13464 11036 13768 11064
rect 11256 10996 11284 11024
rect 10612 10968 11284 10996
rect 12250 10956 12256 11008
rect 12308 10996 12314 11008
rect 13464 10996 13492 11036
rect 12308 10968 13492 10996
rect 12308 10956 12314 10968
rect 13538 10956 13544 11008
rect 13596 10956 13602 11008
rect 13630 10956 13636 11008
rect 13688 10956 13694 11008
rect 13740 11005 13768 11036
rect 13832 11008 13860 11104
rect 14445 11067 14503 11073
rect 14445 11033 14457 11067
rect 14491 11064 14503 11067
rect 14550 11064 14556 11076
rect 14491 11036 14556 11064
rect 14491 11033 14503 11036
rect 14445 11027 14503 11033
rect 14550 11024 14556 11036
rect 14608 11024 14614 11076
rect 14645 11067 14703 11073
rect 14645 11033 14657 11067
rect 14691 11064 14703 11067
rect 14844 11064 14872 11308
rect 15197 11305 15209 11308
rect 15243 11336 15255 11339
rect 16025 11339 16083 11345
rect 16025 11336 16037 11339
rect 15243 11308 16037 11336
rect 15243 11305 15255 11308
rect 15197 11299 15255 11305
rect 16025 11305 16037 11308
rect 16071 11305 16083 11339
rect 19150 11336 19156 11348
rect 16025 11299 16083 11305
rect 18892 11308 19156 11336
rect 14936 11240 15700 11268
rect 14936 11141 14964 11240
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11101 14979 11135
rect 14921 11095 14979 11101
rect 15013 11135 15071 11141
rect 15013 11101 15025 11135
rect 15059 11132 15071 11135
rect 15286 11132 15292 11144
rect 15059 11104 15292 11132
rect 15059 11101 15071 11104
rect 15013 11095 15071 11101
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 15672 11076 15700 11240
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11200 17463 11203
rect 17586 11200 17592 11212
rect 17451 11172 17592 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 17586 11160 17592 11172
rect 17644 11200 17650 11212
rect 18230 11200 18236 11212
rect 17644 11172 18236 11200
rect 17644 11160 17650 11172
rect 18230 11160 18236 11172
rect 18288 11160 18294 11212
rect 18892 11141 18920 11308
rect 19150 11296 19156 11308
rect 19208 11296 19214 11348
rect 19242 11296 19248 11348
rect 19300 11296 19306 11348
rect 19705 11339 19763 11345
rect 19705 11305 19717 11339
rect 19751 11336 19763 11339
rect 19794 11336 19800 11348
rect 19751 11308 19800 11336
rect 19751 11305 19763 11308
rect 19705 11299 19763 11305
rect 19794 11296 19800 11308
rect 19852 11296 19858 11348
rect 20349 11339 20407 11345
rect 20349 11305 20361 11339
rect 20395 11336 20407 11339
rect 20625 11339 20683 11345
rect 20625 11336 20637 11339
rect 20395 11308 20637 11336
rect 20395 11305 20407 11308
rect 20349 11299 20407 11305
rect 20625 11305 20637 11308
rect 20671 11305 20683 11339
rect 20625 11299 20683 11305
rect 20809 11339 20867 11345
rect 20809 11305 20821 11339
rect 20855 11336 20867 11339
rect 21266 11336 21272 11348
rect 20855 11308 21272 11336
rect 20855 11305 20867 11308
rect 20809 11299 20867 11305
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 21358 11296 21364 11348
rect 21416 11296 21422 11348
rect 19061 11271 19119 11277
rect 19061 11237 19073 11271
rect 19107 11268 19119 11271
rect 19334 11268 19340 11280
rect 19107 11240 19340 11268
rect 19107 11237 19119 11240
rect 19061 11231 19119 11237
rect 19334 11228 19340 11240
rect 19392 11228 19398 11280
rect 19886 11228 19892 11280
rect 19944 11228 19950 11280
rect 21376 11268 21404 11296
rect 20180 11240 21404 11268
rect 19797 11203 19855 11209
rect 19797 11200 19809 11203
rect 19444 11172 19809 11200
rect 19444 11141 19472 11172
rect 19797 11169 19809 11172
rect 19843 11200 19855 11203
rect 19904 11200 19932 11228
rect 20180 11200 20208 11240
rect 19843 11172 19932 11200
rect 20088 11172 20208 11200
rect 19843 11169 19855 11172
rect 19797 11163 19855 11169
rect 20088 11141 20116 11172
rect 20622 11160 20628 11212
rect 20680 11160 20686 11212
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11132 19579 11135
rect 20073 11135 20131 11141
rect 20073 11132 20085 11135
rect 19567 11104 20085 11132
rect 19567 11101 19579 11104
rect 19521 11095 19579 11101
rect 20073 11101 20085 11104
rect 20119 11101 20131 11135
rect 20073 11095 20131 11101
rect 20165 11135 20223 11141
rect 20165 11101 20177 11135
rect 20211 11132 20223 11135
rect 20640 11132 20668 11160
rect 20211 11104 20668 11132
rect 20211 11101 20223 11104
rect 20165 11095 20223 11101
rect 14691 11036 14872 11064
rect 15197 11067 15255 11073
rect 14691 11033 14703 11036
rect 14645 11027 14703 11033
rect 15197 11033 15209 11067
rect 15243 11064 15255 11067
rect 15378 11064 15384 11076
rect 15243 11036 15384 11064
rect 15243 11033 15255 11036
rect 15197 11027 15255 11033
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 15654 11024 15660 11076
rect 15712 11064 15718 11076
rect 15712 11036 16068 11064
rect 15712 11024 15718 11036
rect 13725 10999 13783 11005
rect 13725 10965 13737 10999
rect 13771 10965 13783 10999
rect 13725 10959 13783 10965
rect 13814 10956 13820 11008
rect 13872 10956 13878 11008
rect 15930 10956 15936 11008
rect 15988 10956 15994 11008
rect 16040 10996 16068 11036
rect 16850 11024 16856 11076
rect 16908 11064 16914 11076
rect 17138 11067 17196 11073
rect 17138 11064 17150 11067
rect 16908 11036 17150 11064
rect 16908 11024 16914 11036
rect 17138 11033 17150 11036
rect 17184 11033 17196 11067
rect 17138 11027 17196 11033
rect 19705 11067 19763 11073
rect 19705 11033 19717 11067
rect 19751 11064 19763 11067
rect 20180 11064 20208 11095
rect 19751 11036 20208 11064
rect 20441 11067 20499 11073
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 20441 11033 20453 11067
rect 20487 11064 20499 11067
rect 20530 11064 20536 11076
rect 20487 11036 20536 11064
rect 20487 11033 20499 11036
rect 20441 11027 20499 11033
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 20622 11024 20628 11076
rect 20680 11073 20686 11076
rect 20680 11067 20699 11073
rect 20687 11033 20699 11067
rect 20680 11027 20699 11033
rect 20680 11024 20686 11027
rect 17218 10996 17224 11008
rect 16040 10968 17224 10996
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 19981 10999 20039 11005
rect 19981 10996 19993 10999
rect 19852 10968 19993 10996
rect 19852 10956 19858 10968
rect 19981 10965 19993 10968
rect 20027 10965 20039 10999
rect 19981 10959 20039 10965
rect 1104 10906 22264 10928
rect 1104 10854 4255 10906
rect 4307 10854 4319 10906
rect 4371 10854 4383 10906
rect 4435 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 9545 10906
rect 9597 10854 9609 10906
rect 9661 10854 9673 10906
rect 9725 10854 9737 10906
rect 9789 10854 9801 10906
rect 9853 10854 14835 10906
rect 14887 10854 14899 10906
rect 14951 10854 14963 10906
rect 15015 10854 15027 10906
rect 15079 10854 15091 10906
rect 15143 10854 20125 10906
rect 20177 10854 20189 10906
rect 20241 10854 20253 10906
rect 20305 10854 20317 10906
rect 20369 10854 20381 10906
rect 20433 10854 22264 10906
rect 1104 10832 22264 10854
rect 2406 10752 2412 10804
rect 2464 10752 2470 10804
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3329 10795 3387 10801
rect 3329 10792 3341 10795
rect 2832 10764 3341 10792
rect 2832 10752 2838 10764
rect 3329 10761 3341 10764
rect 3375 10761 3387 10795
rect 3329 10755 3387 10761
rect 6181 10795 6239 10801
rect 6181 10761 6193 10795
rect 6227 10792 6239 10795
rect 6362 10792 6368 10804
rect 6227 10764 6368 10792
rect 6227 10761 6239 10764
rect 6181 10755 6239 10761
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 7009 10795 7067 10801
rect 7009 10761 7021 10795
rect 7055 10792 7067 10795
rect 7098 10792 7104 10804
rect 7055 10764 7104 10792
rect 7055 10761 7067 10764
rect 7009 10755 7067 10761
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 7282 10752 7288 10804
rect 7340 10752 7346 10804
rect 7742 10752 7748 10804
rect 7800 10752 7806 10804
rect 8018 10752 8024 10804
rect 8076 10752 8082 10804
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10192 10764 10272 10792
rect 10192 10752 10198 10764
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2424 10656 2452 10752
rect 5068 10727 5126 10733
rect 5068 10693 5080 10727
rect 5114 10724 5126 10727
rect 5994 10724 6000 10736
rect 5114 10696 6000 10724
rect 5114 10693 5126 10696
rect 5068 10687 5126 10693
rect 5994 10684 6000 10696
rect 6052 10684 6058 10736
rect 6380 10724 6408 10752
rect 7300 10724 7328 10752
rect 10244 10733 10272 10764
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11388 10764 11529 10792
rect 11388 10752 11394 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 12802 10752 12808 10804
rect 12860 10752 12866 10804
rect 14550 10752 14556 10804
rect 14608 10792 14614 10804
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 14608 10764 15301 10792
rect 14608 10752 14614 10764
rect 15289 10761 15301 10764
rect 15335 10761 15347 10795
rect 15289 10755 15347 10761
rect 15930 10752 15936 10804
rect 15988 10752 15994 10804
rect 16482 10752 16488 10804
rect 16540 10752 16546 10804
rect 16853 10795 16911 10801
rect 16853 10761 16865 10795
rect 16899 10761 16911 10795
rect 16853 10755 16911 10761
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17218 10792 17224 10804
rect 16991 10764 17224 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 10220 10727 10278 10733
rect 6380 10696 6868 10724
rect 7300 10696 7880 10724
rect 2363 10628 2452 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 3878 10656 3884 10668
rect 3384 10628 3884 10656
rect 3384 10616 3390 10628
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4672 10628 4813 10656
rect 4672 10616 4678 10628
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 6546 10616 6552 10668
rect 6604 10616 6610 10668
rect 6840 10665 6868 10696
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 7006 10616 7012 10668
rect 7064 10656 7070 10668
rect 7852 10665 7880 10696
rect 10220 10693 10232 10727
rect 10266 10693 10278 10727
rect 10220 10687 10278 10693
rect 11606 10684 11612 10736
rect 11664 10684 11670 10736
rect 15427 10693 15485 10699
rect 7101 10659 7159 10665
rect 7101 10656 7113 10659
rect 7064 10628 7113 10656
rect 7064 10616 7070 10628
rect 7101 10625 7113 10628
rect 7147 10625 7159 10659
rect 7101 10619 7159 10625
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 7561 10659 7619 10665
rect 7561 10656 7573 10659
rect 7515 10628 7573 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7561 10625 7573 10628
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10625 7895 10659
rect 11624 10656 11652 10684
rect 15427 10668 15439 10693
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11624 10628 11713 10656
rect 7837 10619 7895 10625
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 2593 10591 2651 10597
rect 2593 10588 2605 10591
rect 2547 10560 2605 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 2593 10557 2605 10560
rect 2639 10557 2651 10591
rect 2593 10551 2651 10557
rect 2958 10548 2964 10600
rect 3016 10588 3022 10600
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 3016 10560 3157 10588
rect 3016 10548 3022 10560
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 3145 10551 3203 10557
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 5960 10560 6653 10588
rect 5960 10548 5966 10560
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 6822 10520 6828 10532
rect 5736 10492 6828 10520
rect 5736 10464 5764 10492
rect 6822 10480 6828 10492
rect 6880 10520 6886 10532
rect 7300 10520 7328 10619
rect 11790 10616 11796 10668
rect 11848 10616 11854 10668
rect 12618 10616 12624 10668
rect 12676 10616 12682 10668
rect 13814 10616 13820 10668
rect 13872 10616 13878 10668
rect 14084 10659 14142 10665
rect 14084 10625 14096 10659
rect 14130 10656 14142 10659
rect 14826 10656 14832 10668
rect 14130 10628 14832 10656
rect 14130 10625 14142 10628
rect 14084 10619 14142 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 15378 10616 15384 10668
rect 15436 10659 15439 10668
rect 15473 10690 15485 10693
rect 15473 10659 15500 10690
rect 15654 10684 15660 10736
rect 15712 10684 15718 10736
rect 15948 10724 15976 10752
rect 15948 10696 16068 10724
rect 15436 10656 15500 10659
rect 15436 10628 15516 10656
rect 15436 10616 15442 10628
rect 9950 10548 9956 10600
rect 10008 10548 10014 10600
rect 13446 10548 13452 10600
rect 13504 10588 13510 10600
rect 13630 10588 13636 10600
rect 13504 10560 13636 10588
rect 13504 10548 13510 10560
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 15488 10588 15516 10628
rect 15930 10616 15936 10668
rect 15988 10616 15994 10668
rect 16040 10665 16068 10696
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10625 16083 10659
rect 16025 10619 16083 10625
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10656 16359 10659
rect 16500 10656 16528 10752
rect 16868 10724 16896 10755
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 18058 10727 18116 10733
rect 18058 10724 18070 10727
rect 16868 10696 18070 10724
rect 18058 10693 18070 10696
rect 18104 10693 18116 10727
rect 18058 10687 18116 10693
rect 19334 10684 19340 10736
rect 19392 10724 19398 10736
rect 19766 10727 19824 10733
rect 19766 10724 19778 10727
rect 19392 10696 19778 10724
rect 19392 10684 19398 10696
rect 19766 10693 19778 10696
rect 19812 10693 19824 10727
rect 19766 10687 19824 10693
rect 16347 10628 16528 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 16666 10616 16672 10668
rect 16724 10616 16730 10668
rect 18230 10616 18236 10668
rect 18288 10656 18294 10668
rect 18325 10659 18383 10665
rect 18325 10656 18337 10659
rect 18288 10628 18337 10656
rect 18288 10616 18294 10628
rect 18325 10625 18337 10628
rect 18371 10656 18383 10659
rect 19521 10659 19579 10665
rect 19521 10656 19533 10659
rect 18371 10628 19533 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 19521 10625 19533 10628
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 16482 10588 16488 10600
rect 15488 10560 16488 10588
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 20993 10591 21051 10597
rect 20993 10557 21005 10591
rect 21039 10557 21051 10591
rect 20993 10551 21051 10557
rect 6880 10492 7328 10520
rect 11333 10523 11391 10529
rect 6880 10480 6886 10492
rect 11333 10489 11345 10523
rect 11379 10520 11391 10523
rect 12250 10520 12256 10532
rect 11379 10492 12256 10520
rect 11379 10489 11391 10492
rect 11333 10483 11391 10489
rect 12250 10480 12256 10492
rect 12308 10480 12314 10532
rect 21008 10464 21036 10551
rect 1946 10412 1952 10464
rect 2004 10452 2010 10464
rect 2133 10455 2191 10461
rect 2133 10452 2145 10455
rect 2004 10424 2145 10452
rect 2004 10412 2010 10424
rect 2133 10421 2145 10424
rect 2179 10421 2191 10455
rect 2133 10415 2191 10421
rect 5718 10412 5724 10464
rect 5776 10412 5782 10464
rect 6638 10412 6644 10464
rect 6696 10412 6702 10464
rect 12066 10412 12072 10464
rect 12124 10412 12130 10464
rect 15197 10455 15255 10461
rect 15197 10421 15209 10455
rect 15243 10452 15255 10455
rect 15286 10452 15292 10464
rect 15243 10424 15292 10452
rect 15243 10421 15255 10424
rect 15197 10415 15255 10421
rect 15286 10412 15292 10424
rect 15344 10452 15350 10464
rect 15473 10455 15531 10461
rect 15473 10452 15485 10455
rect 15344 10424 15485 10452
rect 15344 10412 15350 10424
rect 15473 10421 15485 10424
rect 15519 10421 15531 10455
rect 15473 10415 15531 10421
rect 15746 10412 15752 10464
rect 15804 10412 15810 10464
rect 16485 10455 16543 10461
rect 16485 10421 16497 10455
rect 16531 10452 16543 10455
rect 16850 10452 16856 10464
rect 16531 10424 16856 10452
rect 16531 10421 16543 10424
rect 16485 10415 16543 10421
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 20901 10455 20959 10461
rect 20901 10421 20913 10455
rect 20947 10452 20959 10455
rect 20990 10452 20996 10464
rect 20947 10424 20996 10452
rect 20947 10421 20959 10424
rect 20901 10415 20959 10421
rect 20990 10412 20996 10424
rect 21048 10412 21054 10464
rect 21634 10412 21640 10464
rect 21692 10412 21698 10464
rect 1104 10362 22264 10384
rect 1104 10310 3595 10362
rect 3647 10310 3659 10362
rect 3711 10310 3723 10362
rect 3775 10310 3787 10362
rect 3839 10310 3851 10362
rect 3903 10310 8885 10362
rect 8937 10310 8949 10362
rect 9001 10310 9013 10362
rect 9065 10310 9077 10362
rect 9129 10310 9141 10362
rect 9193 10310 14175 10362
rect 14227 10310 14239 10362
rect 14291 10310 14303 10362
rect 14355 10310 14367 10362
rect 14419 10310 14431 10362
rect 14483 10310 19465 10362
rect 19517 10310 19529 10362
rect 19581 10310 19593 10362
rect 19645 10310 19657 10362
rect 19709 10310 19721 10362
rect 19773 10310 22264 10362
rect 1104 10288 22264 10310
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 3513 10251 3571 10257
rect 3513 10248 3525 10251
rect 3384 10220 3525 10248
rect 3384 10208 3390 10220
rect 3513 10217 3525 10220
rect 3559 10217 3571 10251
rect 3513 10211 3571 10217
rect 4985 10251 5043 10257
rect 4985 10217 4997 10251
rect 5031 10248 5043 10251
rect 5258 10248 5264 10260
rect 5031 10220 5264 10248
rect 5031 10217 5043 10220
rect 4985 10211 5043 10217
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 6549 10251 6607 10257
rect 6549 10248 6561 10251
rect 6012 10220 6561 10248
rect 1578 10072 1584 10124
rect 1636 10112 1642 10124
rect 2133 10115 2191 10121
rect 2133 10112 2145 10115
rect 1636 10084 2145 10112
rect 1636 10072 1642 10084
rect 2133 10081 2145 10084
rect 2179 10081 2191 10115
rect 2133 10075 2191 10081
rect 5902 10072 5908 10124
rect 5960 10112 5966 10124
rect 6012 10121 6040 10220
rect 6549 10217 6561 10220
rect 6595 10217 6607 10251
rect 6549 10211 6607 10217
rect 6730 10208 6736 10260
rect 6788 10208 6794 10260
rect 12066 10208 12072 10260
rect 12124 10208 12130 10260
rect 12526 10208 12532 10260
rect 12584 10208 12590 10260
rect 12894 10208 12900 10260
rect 12952 10208 12958 10260
rect 13357 10251 13415 10257
rect 13357 10217 13369 10251
rect 13403 10248 13415 10251
rect 13630 10248 13636 10260
rect 13403 10220 13636 10248
rect 13403 10217 13415 10220
rect 13357 10211 13415 10217
rect 13630 10208 13636 10220
rect 13688 10248 13694 10260
rect 13688 10220 14688 10248
rect 13688 10208 13694 10220
rect 5997 10115 6055 10121
rect 5997 10112 6009 10115
rect 5960 10084 6009 10112
rect 5960 10072 5966 10084
rect 5997 10081 6009 10084
rect 6043 10081 6055 10115
rect 12084 10112 12112 10208
rect 12912 10180 12940 10208
rect 13541 10183 13599 10189
rect 13541 10180 13553 10183
rect 12912 10152 13553 10180
rect 13541 10149 13553 10152
rect 13587 10149 13599 10183
rect 13541 10143 13599 10149
rect 14660 10121 14688 10220
rect 14826 10208 14832 10260
rect 14884 10208 14890 10260
rect 15746 10248 15752 10260
rect 15212 10220 15752 10248
rect 12161 10115 12219 10121
rect 12161 10112 12173 10115
rect 12084 10084 12173 10112
rect 5997 10075 6055 10081
rect 12161 10081 12173 10084
rect 12207 10081 12219 10115
rect 12161 10075 12219 10081
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10112 13323 10115
rect 14645 10115 14703 10121
rect 13311 10084 13584 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 13556 10056 13584 10084
rect 14645 10081 14657 10115
rect 14691 10081 14703 10115
rect 14645 10075 14703 10081
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 1946 10044 1952 10056
rect 1903 10016 1952 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10013 5227 10047
rect 5169 10007 5227 10013
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10044 5411 10047
rect 5445 10047 5503 10053
rect 5445 10044 5457 10047
rect 5399 10016 5457 10044
rect 5399 10013 5411 10016
rect 5353 10007 5411 10013
rect 5445 10013 5457 10016
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 2378 9979 2436 9985
rect 2378 9976 2390 9979
rect 2056 9948 2390 9976
rect 2056 9917 2084 9948
rect 2378 9945 2390 9948
rect 2424 9945 2436 9979
rect 5184 9976 5212 10007
rect 5718 10004 5724 10056
rect 5776 10004 5782 10056
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 10042 10044 10048 10056
rect 9447 10016 10048 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 5736 9976 5764 10004
rect 5184 9948 5764 9976
rect 2378 9939 2436 9945
rect 6362 9936 6368 9988
rect 6420 9936 6426 9988
rect 6546 9936 6552 9988
rect 6604 9985 6610 9988
rect 6604 9979 6623 9985
rect 6611 9945 6623 9979
rect 9232 9976 9260 10007
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 10318 10004 10324 10056
rect 10376 10004 10382 10056
rect 11606 10004 11612 10056
rect 11664 10044 11670 10056
rect 12342 10044 12348 10056
rect 11664 10016 12348 10044
rect 11664 10004 11670 10016
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 13357 10047 13415 10053
rect 13357 10044 13369 10047
rect 12676 10016 13369 10044
rect 12676 10004 12682 10016
rect 13357 10013 13369 10016
rect 13403 10013 13415 10047
rect 13357 10007 13415 10013
rect 13538 10004 13544 10056
rect 13596 10004 13602 10056
rect 14366 10004 14372 10056
rect 14424 10044 14430 10056
rect 15212 10053 15240 10220
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 20530 10208 20536 10260
rect 20588 10248 20594 10260
rect 20625 10251 20683 10257
rect 20625 10248 20637 10251
rect 20588 10220 20637 10248
rect 20588 10208 20594 10220
rect 20625 10217 20637 10220
rect 20671 10217 20683 10251
rect 20625 10211 20683 10217
rect 16482 10140 16488 10192
rect 16540 10180 16546 10192
rect 16853 10183 16911 10189
rect 16853 10180 16865 10183
rect 16540 10152 16865 10180
rect 16540 10140 16546 10152
rect 16853 10149 16865 10152
rect 16899 10149 16911 10183
rect 20640 10180 20668 10211
rect 20714 10208 20720 10260
rect 20772 10208 20778 10260
rect 20901 10251 20959 10257
rect 20901 10217 20913 10251
rect 20947 10217 20959 10251
rect 20901 10211 20959 10217
rect 20916 10180 20944 10211
rect 21634 10208 21640 10260
rect 21692 10208 21698 10260
rect 20640 10152 20944 10180
rect 16853 10143 16911 10149
rect 16868 10112 16896 10143
rect 21652 10121 21680 10208
rect 17681 10115 17739 10121
rect 17681 10112 17693 10115
rect 16868 10084 17693 10112
rect 17681 10081 17693 10084
rect 17727 10081 17739 10115
rect 21637 10115 21695 10121
rect 17681 10075 17739 10081
rect 20732 10084 21496 10112
rect 20732 10056 20760 10084
rect 15013 10047 15071 10053
rect 15013 10044 15025 10047
rect 14424 10016 15025 10044
rect 14424 10004 14430 10016
rect 15013 10013 15025 10016
rect 15059 10013 15071 10047
rect 15013 10007 15071 10013
rect 15197 10047 15255 10053
rect 15197 10013 15209 10047
rect 15243 10013 15255 10047
rect 15197 10007 15255 10013
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 15436 10016 15485 10044
rect 15436 10004 15442 10016
rect 15473 10013 15485 10016
rect 15519 10013 15531 10047
rect 15473 10007 15531 10013
rect 19058 10004 19064 10056
rect 19116 10004 19122 10056
rect 19245 10047 19303 10053
rect 19245 10013 19257 10047
rect 19291 10044 19303 10047
rect 20530 10044 20536 10056
rect 19291 10016 20536 10044
rect 19291 10013 19303 10016
rect 19245 10007 19303 10013
rect 20530 10004 20536 10016
rect 20588 10004 20594 10056
rect 20714 10004 20720 10056
rect 20772 10004 20778 10056
rect 20898 10004 20904 10056
rect 20956 10004 20962 10056
rect 20990 10004 20996 10056
rect 21048 10004 21054 10056
rect 21468 10053 21496 10084
rect 21637 10081 21649 10115
rect 21683 10081 21695 10115
rect 21637 10075 21695 10081
rect 21453 10047 21511 10053
rect 21453 10013 21465 10047
rect 21499 10013 21511 10047
rect 21453 10007 21511 10013
rect 10336 9976 10364 10004
rect 9232 9948 10364 9976
rect 6604 9939 6623 9945
rect 6604 9936 6610 9939
rect 12250 9936 12256 9988
rect 12308 9976 12314 9988
rect 13081 9979 13139 9985
rect 13081 9976 13093 9979
rect 12308 9948 13093 9976
rect 12308 9936 12314 9948
rect 13081 9945 13093 9948
rect 13127 9945 13139 9979
rect 15718 9979 15776 9985
rect 15718 9976 15730 9979
rect 13081 9939 13139 9945
rect 15396 9948 15730 9976
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9877 2099 9911
rect 2041 9871 2099 9877
rect 9306 9868 9312 9920
rect 9364 9868 9370 9920
rect 14090 9868 14096 9920
rect 14148 9868 14154 9920
rect 15396 9917 15424 9948
rect 15718 9945 15730 9948
rect 15764 9945 15776 9979
rect 15718 9939 15776 9945
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 19490 9979 19548 9985
rect 19490 9976 19502 9979
rect 19392 9948 19502 9976
rect 19392 9936 19398 9948
rect 19490 9945 19502 9948
rect 19536 9945 19548 9979
rect 19490 9939 19548 9945
rect 21082 9936 21088 9988
rect 21140 9976 21146 9988
rect 21177 9979 21235 9985
rect 21177 9976 21189 9979
rect 21140 9948 21189 9976
rect 21140 9936 21146 9948
rect 21177 9945 21189 9948
rect 21223 9945 21235 9979
rect 21177 9939 21235 9945
rect 15381 9911 15439 9917
rect 15381 9877 15393 9911
rect 15427 9877 15439 9911
rect 15381 9871 15439 9877
rect 17129 9911 17187 9917
rect 17129 9877 17141 9911
rect 17175 9908 17187 9911
rect 17218 9908 17224 9920
rect 17175 9880 17224 9908
rect 17175 9877 17187 9880
rect 17129 9871 17187 9877
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 18414 9868 18420 9920
rect 18472 9868 18478 9920
rect 21266 9868 21272 9920
rect 21324 9868 21330 9920
rect 1104 9818 22264 9840
rect 1104 9766 4255 9818
rect 4307 9766 4319 9818
rect 4371 9766 4383 9818
rect 4435 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 9545 9818
rect 9597 9766 9609 9818
rect 9661 9766 9673 9818
rect 9725 9766 9737 9818
rect 9789 9766 9801 9818
rect 9853 9766 14835 9818
rect 14887 9766 14899 9818
rect 14951 9766 14963 9818
rect 15015 9766 15027 9818
rect 15079 9766 15091 9818
rect 15143 9766 20125 9818
rect 20177 9766 20189 9818
rect 20241 9766 20253 9818
rect 20305 9766 20317 9818
rect 20369 9766 20381 9818
rect 20433 9766 22264 9818
rect 1104 9744 22264 9766
rect 2958 9664 2964 9716
rect 3016 9664 3022 9716
rect 9861 9707 9919 9713
rect 5368 9676 7880 9704
rect 3142 9596 3148 9648
rect 3200 9636 3206 9648
rect 4062 9636 4068 9648
rect 3200 9608 4068 9636
rect 3200 9596 3206 9608
rect 1578 9528 1584 9580
rect 1636 9528 1642 9580
rect 1848 9571 1906 9577
rect 1848 9537 1860 9571
rect 1894 9568 1906 9571
rect 2222 9568 2228 9580
rect 1894 9540 2228 9568
rect 1894 9537 1906 9540
rect 1848 9531 1906 9537
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 3988 9577 4016 9608
rect 4062 9596 4068 9608
rect 4120 9636 4126 9648
rect 5368 9636 5396 9676
rect 7852 9636 7880 9676
rect 9861 9673 9873 9707
rect 9907 9704 9919 9707
rect 10042 9704 10048 9716
rect 9907 9676 10048 9704
rect 9907 9673 9919 9676
rect 9861 9667 9919 9673
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 12342 9664 12348 9716
rect 12400 9704 12406 9716
rect 16022 9704 16028 9716
rect 12400 9676 16028 9704
rect 12400 9664 12406 9676
rect 8021 9639 8079 9645
rect 8021 9636 8033 9639
rect 4120 9608 5396 9636
rect 5460 9608 7788 9636
rect 7852 9608 8033 9636
rect 4120 9596 4126 9608
rect 5460 9577 5488 9608
rect 7760 9580 7788 9608
rect 8021 9605 8033 9608
rect 8067 9636 8079 9639
rect 8067 9608 8432 9636
rect 8067 9605 8079 9608
rect 8021 9599 8079 9605
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9537 5503 9571
rect 5445 9531 5503 9537
rect 4172 9500 4200 9531
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 5813 9571 5871 9577
rect 5592 9566 5764 9568
rect 5813 9566 5825 9571
rect 5592 9540 5825 9566
rect 5592 9528 5598 9540
rect 5736 9538 5825 9540
rect 5813 9537 5825 9538
rect 5859 9537 5871 9571
rect 5813 9531 5871 9537
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9537 5963 9571
rect 5905 9531 5963 9537
rect 6089 9571 6147 9577
rect 6089 9537 6101 9571
rect 6135 9568 6147 9571
rect 6362 9568 6368 9580
rect 6135 9540 6368 9568
rect 6135 9537 6147 9540
rect 6089 9531 6147 9537
rect 4338 9500 4344 9512
rect 4172 9472 4344 9500
rect 4338 9460 4344 9472
rect 4396 9500 4402 9512
rect 5721 9503 5779 9509
rect 5721 9500 5733 9503
rect 4396 9472 5733 9500
rect 4396 9460 4402 9472
rect 5721 9469 5733 9472
rect 5767 9469 5779 9503
rect 5721 9463 5779 9469
rect 5920 9432 5948 9531
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7300 9444 7328 9531
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9537 8263 9571
rect 8205 9531 8263 9537
rect 8220 9500 8248 9531
rect 8294 9528 8300 9580
rect 8352 9528 8358 9580
rect 8404 9568 8432 9608
rect 9306 9596 9312 9648
rect 9364 9636 9370 9648
rect 9502 9639 9560 9645
rect 9502 9636 9514 9639
rect 9364 9608 9514 9636
rect 9364 9596 9370 9608
rect 9502 9605 9514 9608
rect 9548 9605 9560 9639
rect 10778 9636 10784 9648
rect 9502 9599 9560 9605
rect 9600 9608 10784 9636
rect 9600 9568 9628 9608
rect 10778 9596 10784 9608
rect 10836 9596 10842 9648
rect 8404 9540 9628 9568
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 10410 9568 10416 9580
rect 10336 9540 10416 9568
rect 8662 9500 8668 9512
rect 8220 9472 8668 9500
rect 8662 9460 8668 9472
rect 8720 9460 8726 9512
rect 9769 9503 9827 9509
rect 9769 9469 9781 9503
rect 9815 9500 9827 9503
rect 9950 9500 9956 9512
rect 9815 9472 9956 9500
rect 9815 9469 9827 9472
rect 9769 9463 9827 9469
rect 5092 9404 5948 9432
rect 5092 9376 5120 9404
rect 7282 9392 7288 9444
rect 7340 9392 7346 9444
rect 8220 9404 8892 9432
rect 8220 9376 8248 9404
rect 3970 9324 3976 9376
rect 4028 9324 4034 9376
rect 5074 9324 5080 9376
rect 5132 9324 5138 9376
rect 5258 9324 5264 9376
rect 5316 9324 5322 9376
rect 5626 9324 5632 9376
rect 5684 9324 5690 9376
rect 6086 9324 6092 9376
rect 6144 9324 6150 9376
rect 7193 9367 7251 9373
rect 7193 9333 7205 9367
rect 7239 9364 7251 9367
rect 7374 9364 7380 9376
rect 7239 9336 7380 9364
rect 7239 9333 7251 9336
rect 7193 9327 7251 9333
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 8021 9367 8079 9373
rect 8021 9333 8033 9367
rect 8067 9364 8079 9367
rect 8110 9364 8116 9376
rect 8067 9336 8116 9364
rect 8067 9333 8079 9336
rect 8021 9327 8079 9333
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 8202 9324 8208 9376
rect 8260 9324 8266 9376
rect 8386 9324 8392 9376
rect 8444 9324 8450 9376
rect 8864 9364 8892 9404
rect 9784 9364 9812 9463
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 10042 9460 10048 9512
rect 10100 9500 10106 9512
rect 10100 9472 10145 9500
rect 10100 9460 10106 9472
rect 10226 9460 10232 9512
rect 10284 9460 10290 9512
rect 10336 9509 10364 9540
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 10594 9528 10600 9580
rect 10652 9568 10658 9580
rect 11609 9571 11667 9577
rect 11609 9568 11621 9571
rect 10652 9540 11621 9568
rect 10652 9528 10658 9540
rect 11609 9537 11621 9540
rect 11655 9537 11667 9571
rect 11609 9531 11667 9537
rect 11790 9528 11796 9580
rect 11848 9528 11854 9580
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13648 9568 13676 9676
rect 14568 9648 14596 9676
rect 16022 9664 16028 9676
rect 16080 9704 16086 9716
rect 16080 9676 16620 9704
rect 16080 9664 16086 9676
rect 13725 9639 13783 9645
rect 13725 9605 13737 9639
rect 13771 9636 13783 9639
rect 14366 9636 14372 9648
rect 13771 9608 14372 9636
rect 13771 9605 13783 9608
rect 13725 9599 13783 9605
rect 14366 9596 14372 9608
rect 14424 9596 14430 9648
rect 14550 9596 14556 9648
rect 14608 9596 14614 9648
rect 13587 9540 13676 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 14090 9528 14096 9580
rect 14148 9528 14154 9580
rect 16592 9568 16620 9676
rect 16666 9664 16672 9716
rect 16724 9704 16730 9716
rect 16945 9707 17003 9713
rect 16945 9704 16957 9707
rect 16724 9676 16957 9704
rect 16724 9664 16730 9676
rect 16945 9673 16957 9676
rect 16991 9673 17003 9707
rect 16945 9667 17003 9673
rect 19058 9664 19064 9716
rect 19116 9704 19122 9716
rect 19153 9707 19211 9713
rect 19153 9704 19165 9707
rect 19116 9676 19165 9704
rect 19116 9664 19122 9676
rect 19153 9673 19165 9676
rect 19199 9673 19211 9707
rect 19153 9667 19211 9673
rect 20793 9707 20851 9713
rect 20793 9673 20805 9707
rect 20839 9704 20851 9707
rect 21082 9704 21088 9716
rect 20839 9676 21088 9704
rect 20839 9673 20851 9676
rect 20793 9667 20851 9673
rect 19168 9636 19196 9667
rect 21082 9664 21088 9676
rect 21140 9664 21146 9716
rect 21266 9664 21272 9716
rect 21324 9664 21330 9716
rect 20898 9636 20904 9648
rect 19168 9608 20904 9636
rect 20898 9596 20904 9608
rect 20956 9636 20962 9648
rect 20993 9639 21051 9645
rect 20993 9636 21005 9639
rect 20956 9608 21005 9636
rect 20956 9596 20962 9608
rect 20993 9605 21005 9608
rect 21039 9605 21051 9639
rect 20993 9599 21051 9605
rect 17129 9571 17187 9577
rect 17129 9568 17141 9571
rect 16592 9540 17141 9568
rect 17129 9537 17141 9540
rect 17175 9537 17187 9571
rect 17129 9531 17187 9537
rect 18414 9528 18420 9580
rect 18472 9528 18478 9580
rect 18598 9528 18604 9580
rect 18656 9528 18662 9580
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9568 18843 9571
rect 18877 9571 18935 9577
rect 18877 9568 18889 9571
rect 18831 9540 18889 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 18877 9537 18889 9540
rect 18923 9537 18935 9571
rect 18877 9531 18935 9537
rect 20277 9571 20335 9577
rect 20277 9537 20289 9571
rect 20323 9568 20335 9571
rect 20438 9568 20444 9580
rect 20323 9540 20444 9568
rect 20323 9537 20335 9540
rect 20277 9531 20335 9537
rect 20438 9528 20444 9540
rect 20496 9528 20502 9580
rect 21284 9577 21312 9664
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9537 21327 9571
rect 21269 9531 21327 9537
rect 10321 9503 10379 9509
rect 10321 9469 10333 9503
rect 10367 9469 10379 9503
rect 11882 9500 11888 9512
rect 10321 9463 10379 9469
rect 10513 9472 11888 9500
rect 10410 9392 10416 9444
rect 10468 9432 10474 9444
rect 10513 9432 10541 9472
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9500 13415 9503
rect 14108 9500 14136 9528
rect 13403 9472 14136 9500
rect 13403 9469 13415 9472
rect 13357 9463 13415 9469
rect 17218 9460 17224 9512
rect 17276 9500 17282 9512
rect 17313 9503 17371 9509
rect 17313 9500 17325 9503
rect 17276 9472 17325 9500
rect 17276 9460 17282 9472
rect 17313 9469 17325 9472
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 20530 9460 20536 9512
rect 20588 9460 20594 9512
rect 10468 9404 10541 9432
rect 19061 9435 19119 9441
rect 10468 9392 10474 9404
rect 19061 9401 19073 9435
rect 19107 9432 19119 9435
rect 19334 9432 19340 9444
rect 19107 9404 19340 9432
rect 19107 9401 19119 9404
rect 19061 9395 19119 9401
rect 19334 9392 19340 9404
rect 19392 9392 19398 9444
rect 20622 9392 20628 9444
rect 20680 9392 20686 9444
rect 8864 9336 9812 9364
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 11793 9367 11851 9373
rect 11793 9364 11805 9367
rect 11664 9336 11805 9364
rect 11664 9324 11670 9336
rect 11793 9333 11805 9336
rect 11839 9333 11851 9367
rect 11793 9327 11851 9333
rect 20809 9367 20867 9373
rect 20809 9333 20821 9367
rect 20855 9364 20867 9367
rect 20990 9364 20996 9376
rect 20855 9336 20996 9364
rect 20855 9333 20867 9336
rect 20809 9327 20867 9333
rect 20990 9324 20996 9336
rect 21048 9324 21054 9376
rect 21082 9324 21088 9376
rect 21140 9324 21146 9376
rect 1104 9274 22264 9296
rect 1104 9222 3595 9274
rect 3647 9222 3659 9274
rect 3711 9222 3723 9274
rect 3775 9222 3787 9274
rect 3839 9222 3851 9274
rect 3903 9222 8885 9274
rect 8937 9222 8949 9274
rect 9001 9222 9013 9274
rect 9065 9222 9077 9274
rect 9129 9222 9141 9274
rect 9193 9222 14175 9274
rect 14227 9222 14239 9274
rect 14291 9222 14303 9274
rect 14355 9222 14367 9274
rect 14419 9222 14431 9274
rect 14483 9222 19465 9274
rect 19517 9222 19529 9274
rect 19581 9222 19593 9274
rect 19645 9222 19657 9274
rect 19709 9222 19721 9274
rect 19773 9222 22264 9274
rect 1104 9200 22264 9222
rect 2222 9120 2228 9172
rect 2280 9120 2286 9172
rect 4062 9120 4068 9172
rect 4120 9120 4126 9172
rect 4338 9120 4344 9172
rect 4396 9120 4402 9172
rect 5626 9120 5632 9172
rect 5684 9160 5690 9172
rect 5905 9163 5963 9169
rect 5905 9160 5917 9163
rect 5684 9132 5917 9160
rect 5684 9120 5690 9132
rect 5905 9129 5917 9132
rect 5951 9129 5963 9163
rect 5905 9123 5963 9129
rect 6086 9120 6092 9172
rect 6144 9120 6150 9172
rect 8110 9120 8116 9172
rect 8168 9120 8174 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8573 9163 8631 9169
rect 8573 9160 8585 9163
rect 8352 9132 8585 9160
rect 8352 9120 8358 9132
rect 8573 9129 8585 9132
rect 8619 9160 8631 9163
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 8619 9132 8953 9160
rect 8619 9129 8631 9132
rect 8573 9123 8631 9129
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 10042 9160 10048 9172
rect 8941 9123 8999 9129
rect 9324 9132 10048 9160
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9061 1639 9095
rect 1581 9055 1639 9061
rect 1596 9024 1624 9055
rect 3973 9027 4031 9033
rect 1596 8996 1992 9024
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1854 8916 1860 8968
rect 1912 8916 1918 8968
rect 1964 8965 1992 8996
rect 3973 8993 3985 9027
rect 4019 9024 4031 9027
rect 4080 9024 4108 9120
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 4019 8996 4108 9024
rect 4264 8996 5181 9024
rect 4019 8993 4031 8996
rect 3973 8987 4031 8993
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8925 2007 8959
rect 1949 8919 2007 8925
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8956 2191 8959
rect 2409 8959 2467 8965
rect 2409 8956 2421 8959
rect 2179 8928 2421 8956
rect 2179 8925 2191 8928
rect 2133 8919 2191 8925
rect 2409 8925 2421 8928
rect 2455 8925 2467 8959
rect 2409 8919 2467 8925
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4264 8965 4292 8996
rect 5169 8993 5181 8996
rect 5215 8993 5227 9027
rect 5169 8987 5227 8993
rect 5534 8984 5540 9036
rect 5592 8984 5598 9036
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 9024 5871 9027
rect 6104 9024 6132 9120
rect 5859 8996 6132 9024
rect 8128 9024 8156 9120
rect 8128 8996 8432 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 4120 8928 4169 8956
rect 4120 8916 4126 8928
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5074 8956 5080 8968
rect 5031 8928 5080 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 5552 8956 5580 8984
rect 6086 8956 6092 8968
rect 5552 8928 6092 8956
rect 6086 8916 6092 8928
rect 6144 8956 6150 8968
rect 6549 8959 6607 8965
rect 6549 8956 6561 8959
rect 6144 8928 6561 8956
rect 6144 8916 6150 8928
rect 6549 8925 6561 8928
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 8113 8959 8171 8965
rect 8113 8925 8125 8959
rect 8159 8956 8171 8959
rect 8202 8956 8208 8968
rect 8159 8928 8208 8956
rect 8159 8925 8171 8928
rect 8113 8919 8171 8925
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 8404 8965 8432 8996
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9324 9024 9352 9132
rect 10042 9120 10048 9132
rect 10100 9160 10106 9172
rect 10410 9160 10416 9172
rect 10100 9132 10416 9160
rect 10100 9120 10106 9132
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 11422 9120 11428 9172
rect 11480 9160 11486 9172
rect 11480 9132 11560 9160
rect 11480 9120 11486 9132
rect 9953 9095 10011 9101
rect 9953 9092 9965 9095
rect 9088 8996 9352 9024
rect 9088 8984 9094 8996
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 8665 8959 8723 8965
rect 8665 8925 8677 8959
rect 8711 8925 8723 8959
rect 8665 8919 8723 8925
rect 7868 8891 7926 8897
rect 7868 8857 7880 8891
rect 7914 8888 7926 8891
rect 7914 8860 8248 8888
rect 7914 8857 7926 8860
rect 7868 8851 7926 8857
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 4249 8823 4307 8829
rect 4249 8820 4261 8823
rect 4212 8792 4261 8820
rect 4212 8780 4218 8792
rect 4249 8789 4261 8792
rect 4295 8789 4307 8823
rect 4249 8783 4307 8789
rect 6733 8823 6791 8829
rect 6733 8789 6745 8823
rect 6779 8820 6791 8823
rect 7282 8820 7288 8832
rect 6779 8792 7288 8820
rect 6779 8789 6791 8792
rect 6733 8783 6791 8789
rect 7282 8780 7288 8792
rect 7340 8820 7346 8832
rect 8018 8820 8024 8832
rect 7340 8792 8024 8820
rect 7340 8780 7346 8792
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8220 8829 8248 8860
rect 8680 8832 8708 8919
rect 9214 8916 9220 8968
rect 9272 8916 9278 8968
rect 9324 8965 9352 8996
rect 9416 9064 9965 9092
rect 9416 8965 9444 9064
rect 9953 9061 9965 9064
rect 9999 9092 10011 9095
rect 10229 9095 10287 9101
rect 10229 9092 10241 9095
rect 9999 9064 10241 9092
rect 9999 9061 10011 9064
rect 9953 9055 10011 9061
rect 10229 9061 10241 9064
rect 10275 9061 10287 9095
rect 10229 9055 10287 9061
rect 10502 9052 10508 9104
rect 10560 9092 10566 9104
rect 11146 9092 11152 9104
rect 10560 9064 11152 9092
rect 10560 9052 10566 9064
rect 11146 9052 11152 9064
rect 11204 9052 11210 9104
rect 11532 9092 11560 9132
rect 11790 9120 11796 9172
rect 11848 9120 11854 9172
rect 11882 9120 11888 9172
rect 11940 9120 11946 9172
rect 13538 9120 13544 9172
rect 13596 9160 13602 9172
rect 14093 9163 14151 9169
rect 14093 9160 14105 9163
rect 13596 9132 14105 9160
rect 13596 9120 13602 9132
rect 14093 9129 14105 9132
rect 14139 9129 14151 9163
rect 14093 9123 14151 9129
rect 20438 9120 20444 9172
rect 20496 9120 20502 9172
rect 21174 9120 21180 9172
rect 21232 9160 21238 9172
rect 21913 9163 21971 9169
rect 21913 9160 21925 9163
rect 21232 9132 21925 9160
rect 21232 9120 21238 9132
rect 21913 9129 21925 9132
rect 21959 9129 21971 9163
rect 21913 9123 21971 9129
rect 11532 9064 12848 9092
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 11238 9024 11244 9036
rect 10468 8996 11244 9024
rect 10468 8984 10474 8996
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 9585 8959 9643 8965
rect 9585 8925 9597 8959
rect 9631 8956 9643 8959
rect 10226 8956 10232 8968
rect 9631 8928 10232 8956
rect 9631 8925 9643 8928
rect 9585 8919 9643 8925
rect 9416 8888 9444 8919
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 11072 8965 11100 8996
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 11330 8984 11336 9036
rect 11388 8984 11394 9036
rect 11422 8984 11428 9036
rect 11480 8984 11486 9036
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 10560 8928 10885 8956
rect 10560 8916 10566 8928
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8925 11115 8959
rect 11057 8919 11115 8925
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8956 11207 8959
rect 11514 8956 11520 8968
rect 11195 8950 11284 8956
rect 11440 8950 11520 8956
rect 11195 8928 11520 8950
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 11256 8922 11468 8928
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 11698 8956 11704 8968
rect 11655 8928 11704 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 12066 8916 12072 8968
rect 12124 8916 12130 8968
rect 12345 8959 12403 8965
rect 12345 8925 12357 8959
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 12529 8959 12587 8965
rect 12529 8925 12541 8959
rect 12575 8956 12587 8959
rect 12710 8956 12716 8968
rect 12575 8928 12716 8956
rect 12575 8925 12587 8928
rect 12529 8919 12587 8925
rect 9140 8860 9444 8888
rect 9140 8832 9168 8860
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 9677 8891 9735 8897
rect 9677 8888 9689 8891
rect 9548 8860 9689 8888
rect 9548 8848 9554 8860
rect 9677 8857 9689 8860
rect 9723 8857 9735 8891
rect 10413 8891 10471 8897
rect 10413 8888 10425 8891
rect 9677 8851 9735 8857
rect 9876 8860 10425 8888
rect 8205 8823 8263 8829
rect 8205 8789 8217 8823
rect 8251 8789 8263 8823
rect 8205 8783 8263 8789
rect 8662 8780 8668 8832
rect 8720 8780 8726 8832
rect 9122 8780 9128 8832
rect 9180 8780 9186 8832
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 9876 8820 9904 8860
rect 10413 8857 10425 8860
rect 10459 8857 10471 8891
rect 10413 8851 10471 8857
rect 10597 8891 10655 8897
rect 10597 8857 10609 8891
rect 10643 8888 10655 8891
rect 12360 8888 12388 8919
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 12820 8965 12848 9064
rect 19978 9052 19984 9104
rect 20036 9052 20042 9104
rect 19996 9024 20024 9052
rect 17236 8996 20024 9024
rect 12805 8959 12863 8965
rect 12805 8925 12817 8959
rect 12851 8956 12863 8959
rect 12851 8928 13492 8956
rect 12851 8925 12863 8928
rect 12805 8919 12863 8925
rect 10643 8860 10824 8888
rect 10643 8857 10655 8860
rect 10597 8851 10655 8857
rect 9364 8792 9904 8820
rect 9364 8780 9370 8792
rect 10134 8780 10140 8832
rect 10192 8780 10198 8832
rect 10686 8780 10692 8832
rect 10744 8780 10750 8832
rect 10796 8820 10824 8860
rect 11440 8860 12388 8888
rect 11054 8820 11060 8832
rect 10796 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8820 11118 8832
rect 11440 8820 11468 8860
rect 13464 8832 13492 8928
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 15473 8959 15531 8965
rect 15473 8956 15485 8959
rect 15436 8928 15485 8956
rect 15436 8916 15442 8928
rect 15473 8925 15485 8928
rect 15519 8925 15531 8959
rect 15473 8919 15531 8925
rect 16114 8916 16120 8968
rect 16172 8916 16178 8968
rect 16850 8916 16856 8968
rect 16908 8956 16914 8968
rect 17236 8965 17264 8996
rect 20530 8984 20536 9036
rect 20588 8984 20594 9036
rect 17221 8959 17279 8965
rect 17221 8956 17233 8959
rect 16908 8928 17233 8956
rect 16908 8916 16914 8928
rect 17221 8925 17233 8928
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 17402 8916 17408 8968
rect 17460 8916 17466 8968
rect 19886 8916 19892 8968
rect 19944 8916 19950 8968
rect 19981 8959 20039 8965
rect 19981 8925 19993 8959
rect 20027 8925 20039 8959
rect 19981 8919 20039 8925
rect 20165 8959 20223 8965
rect 20165 8925 20177 8959
rect 20211 8956 20223 8959
rect 20257 8959 20315 8965
rect 20257 8956 20269 8959
rect 20211 8928 20269 8956
rect 20211 8925 20223 8928
rect 20165 8919 20223 8925
rect 20257 8925 20269 8928
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 20800 8959 20858 8965
rect 20800 8925 20812 8959
rect 20846 8956 20858 8959
rect 21082 8956 21088 8968
rect 20846 8928 21088 8956
rect 20846 8925 20858 8928
rect 20800 8919 20858 8925
rect 15194 8848 15200 8900
rect 15252 8897 15258 8900
rect 15252 8851 15264 8897
rect 16132 8888 16160 8916
rect 19996 8888 20024 8919
rect 21082 8916 21088 8928
rect 21140 8916 21146 8968
rect 20714 8888 20720 8900
rect 16132 8860 20720 8888
rect 15252 8848 15258 8851
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 11112 8792 11468 8820
rect 11112 8780 11118 8792
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 12713 8823 12771 8829
rect 12713 8820 12725 8823
rect 12400 8792 12725 8820
rect 12400 8780 12406 8792
rect 12713 8789 12725 8792
rect 12759 8789 12771 8823
rect 12713 8783 12771 8789
rect 13446 8780 13452 8832
rect 13504 8780 13510 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 17037 8823 17095 8829
rect 17037 8820 17049 8823
rect 16632 8792 17049 8820
rect 16632 8780 16638 8792
rect 17037 8789 17049 8792
rect 17083 8789 17095 8823
rect 17037 8783 17095 8789
rect 1104 8730 22264 8752
rect 1104 8678 4255 8730
rect 4307 8678 4319 8730
rect 4371 8678 4383 8730
rect 4435 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 9545 8730
rect 9597 8678 9609 8730
rect 9661 8678 9673 8730
rect 9725 8678 9737 8730
rect 9789 8678 9801 8730
rect 9853 8678 14835 8730
rect 14887 8678 14899 8730
rect 14951 8678 14963 8730
rect 15015 8678 15027 8730
rect 15079 8678 15091 8730
rect 15143 8678 20125 8730
rect 20177 8678 20189 8730
rect 20241 8678 20253 8730
rect 20305 8678 20317 8730
rect 20369 8678 20381 8730
rect 20433 8678 22264 8730
rect 1104 8656 22264 8678
rect 3970 8576 3976 8628
rect 4028 8576 4034 8628
rect 5258 8576 5264 8628
rect 5316 8576 5322 8628
rect 6086 8576 6092 8628
rect 6144 8576 6150 8628
rect 6362 8576 6368 8628
rect 6420 8576 6426 8628
rect 9030 8576 9036 8628
rect 9088 8576 9094 8628
rect 9398 8576 9404 8628
rect 9456 8616 9462 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9456 8588 9505 8616
rect 9456 8576 9462 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 9493 8579 9551 8585
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 10008 8588 10057 8616
rect 10008 8576 10014 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10045 8579 10103 8585
rect 10498 8619 10556 8625
rect 10498 8585 10510 8619
rect 10544 8616 10556 8619
rect 10594 8616 10600 8628
rect 10544 8588 10600 8616
rect 10544 8585 10556 8588
rect 10498 8579 10556 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 10686 8576 10692 8628
rect 10744 8576 10750 8628
rect 11330 8576 11336 8628
rect 11388 8576 11394 8628
rect 11698 8616 11704 8628
rect 11440 8588 11704 8616
rect 3412 8551 3470 8557
rect 3412 8517 3424 8551
rect 3458 8548 3470 8551
rect 3988 8548 4016 8576
rect 3458 8520 4016 8548
rect 4976 8551 5034 8557
rect 3458 8517 3470 8520
rect 3412 8511 3470 8517
rect 4976 8517 4988 8551
rect 5022 8548 5034 8551
rect 5276 8548 5304 8576
rect 5022 8520 5304 8548
rect 5022 8517 5034 8520
rect 4976 8511 5034 8517
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 8113 8551 8171 8557
rect 8113 8548 8125 8551
rect 7064 8520 8125 8548
rect 7064 8508 7070 8520
rect 8113 8517 8125 8520
rect 8159 8517 8171 8551
rect 8113 8511 8171 8517
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 1636 8452 3188 8480
rect 1636 8440 1642 8452
rect 3160 8421 3188 8452
rect 7374 8440 7380 8492
rect 7432 8480 7438 8492
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 7432 8452 7573 8480
rect 7432 8440 7438 8452
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7650 8440 7656 8492
rect 7708 8480 7714 8492
rect 8021 8483 8079 8489
rect 8021 8480 8033 8483
rect 7708 8452 8033 8480
rect 7708 8440 7714 8452
rect 8021 8449 8033 8452
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8294 8440 8300 8492
rect 8352 8440 8358 8492
rect 9048 8489 9076 8576
rect 9122 8508 9128 8560
rect 9180 8508 9186 8560
rect 8941 8483 8999 8489
rect 8941 8449 8953 8483
rect 8987 8449 8999 8483
rect 8941 8443 8999 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 3145 8415 3203 8421
rect 3145 8381 3157 8415
rect 3191 8381 3203 8415
rect 3145 8375 3203 8381
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8381 4767 8415
rect 4709 8375 4767 8381
rect 3160 8276 3188 8375
rect 4724 8344 4752 8375
rect 6914 8372 6920 8424
rect 6972 8372 6978 8424
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8412 7527 8415
rect 7834 8412 7840 8424
rect 7515 8384 7840 8412
rect 7515 8381 7527 8384
rect 7469 8375 7527 8381
rect 7834 8372 7840 8384
rect 7892 8372 7898 8424
rect 8662 8412 8668 8424
rect 7944 8384 8668 8412
rect 7944 8353 7972 8384
rect 8662 8372 8668 8384
rect 8720 8412 8726 8424
rect 8956 8412 8984 8443
rect 9214 8440 9220 8492
rect 9272 8440 9278 8492
rect 9416 8489 9444 8576
rect 9858 8508 9864 8560
rect 9916 8548 9922 8560
rect 10229 8551 10287 8557
rect 9916 8520 10180 8548
rect 9916 8508 9922 8520
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 9582 8440 9588 8492
rect 9640 8480 9646 8492
rect 9677 8483 9735 8489
rect 9677 8480 9689 8483
rect 9640 8452 9689 8480
rect 9640 8440 9646 8452
rect 9677 8449 9689 8452
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 9953 8483 10011 8489
rect 9953 8449 9965 8483
rect 9999 8449 10011 8483
rect 10152 8480 10180 8520
rect 10229 8517 10241 8551
rect 10275 8548 10287 8551
rect 10704 8548 10732 8576
rect 10275 8520 10732 8548
rect 10275 8517 10287 8520
rect 10229 8511 10287 8517
rect 10321 8483 10379 8489
rect 10321 8480 10333 8483
rect 10152 8452 10333 8480
rect 9953 8443 10011 8449
rect 10321 8449 10333 8452
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 9861 8415 9919 8421
rect 9861 8412 9873 8415
rect 8720 8384 8984 8412
rect 9508 8384 9873 8412
rect 8720 8372 8726 8384
rect 4080 8316 4752 8344
rect 7929 8347 7987 8353
rect 3510 8276 3516 8288
rect 3160 8248 3516 8276
rect 3510 8236 3516 8248
rect 3568 8276 3574 8288
rect 4080 8276 4108 8316
rect 7929 8313 7941 8347
rect 7975 8313 7987 8347
rect 7929 8307 7987 8313
rect 8386 8304 8392 8356
rect 8444 8304 8450 8356
rect 8478 8304 8484 8356
rect 8536 8304 8542 8356
rect 8757 8347 8815 8353
rect 8757 8313 8769 8347
rect 8803 8344 8815 8347
rect 9398 8344 9404 8356
rect 8803 8316 9404 8344
rect 8803 8313 8815 8316
rect 8757 8307 8815 8313
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 3568 8248 4108 8276
rect 4525 8279 4583 8285
rect 3568 8236 3574 8248
rect 4525 8245 4537 8279
rect 4571 8276 4583 8279
rect 5074 8276 5080 8288
rect 4571 8248 5080 8276
rect 4571 8245 4583 8248
rect 4525 8239 4583 8245
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 8404 8276 8432 8304
rect 9306 8276 9312 8288
rect 8404 8248 9312 8276
rect 9306 8236 9312 8248
rect 9364 8276 9370 8288
rect 9508 8276 9536 8384
rect 9861 8381 9873 8384
rect 9907 8381 9919 8415
rect 9968 8412 9996 8443
rect 10410 8440 10416 8492
rect 10468 8440 10474 8492
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 11440 8480 11468 8588
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 12897 8619 12955 8625
rect 12897 8616 12909 8619
rect 12768 8588 12909 8616
rect 12768 8576 12774 8588
rect 12897 8585 12909 8588
rect 12943 8616 12955 8619
rect 16025 8619 16083 8625
rect 12943 8588 13768 8616
rect 12943 8585 12955 8588
rect 12897 8579 12955 8585
rect 10643 8452 11468 8480
rect 11532 8520 13584 8548
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 10686 8412 10692 8424
rect 9968 8384 10692 8412
rect 9861 8375 9919 8381
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11422 8412 11428 8424
rect 10827 8384 11428 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 11422 8372 11428 8384
rect 11480 8372 11486 8424
rect 11532 8421 11560 8520
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 11773 8483 11831 8489
rect 11773 8480 11785 8483
rect 11664 8452 11785 8480
rect 11664 8440 11670 8452
rect 11773 8449 11785 8452
rect 11819 8449 11831 8483
rect 11773 8443 11831 8449
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8381 11575 8415
rect 13556 8412 13584 8520
rect 13630 8440 13636 8492
rect 13688 8440 13694 8492
rect 13740 8489 13768 8588
rect 16025 8585 16037 8619
rect 16071 8616 16083 8619
rect 16114 8616 16120 8628
rect 16071 8588 16120 8616
rect 16071 8585 16083 8588
rect 16025 8579 16083 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16485 8619 16543 8625
rect 16485 8585 16497 8619
rect 16531 8616 16543 8619
rect 16531 8588 16804 8616
rect 16531 8585 16543 8588
rect 16485 8579 16543 8585
rect 15378 8548 15384 8560
rect 14016 8520 15384 8548
rect 13725 8483 13783 8489
rect 13725 8449 13737 8483
rect 13771 8449 13783 8483
rect 13725 8443 13783 8449
rect 14016 8421 14044 8520
rect 15378 8508 15384 8520
rect 15436 8548 15442 8560
rect 16776 8548 16804 8588
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 18141 8619 18199 8625
rect 18141 8616 18153 8619
rect 17460 8588 18153 8616
rect 17460 8576 17466 8588
rect 18141 8585 18153 8588
rect 18187 8585 18199 8619
rect 18141 8579 18199 8585
rect 19886 8576 19892 8628
rect 19944 8616 19950 8628
rect 20901 8619 20959 8625
rect 20901 8616 20913 8619
rect 19944 8588 20913 8616
rect 19944 8576 19950 8588
rect 20901 8585 20913 8588
rect 20947 8585 20959 8619
rect 20901 8579 20959 8585
rect 16914 8551 16972 8557
rect 16914 8548 16926 8551
rect 15436 8520 16712 8548
rect 16776 8520 16926 8548
rect 15436 8508 15442 8520
rect 14090 8440 14096 8492
rect 14148 8480 14154 8492
rect 14257 8483 14315 8489
rect 14257 8480 14269 8483
rect 14148 8452 14269 8480
rect 14148 8440 14154 8452
rect 14257 8449 14269 8452
rect 14303 8449 14315 8483
rect 14257 8443 14315 8449
rect 15838 8440 15844 8492
rect 15896 8440 15902 8492
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 16574 8480 16580 8492
rect 16347 8452 16580 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 16684 8489 16712 8520
rect 16914 8517 16926 8520
rect 16960 8517 16972 8551
rect 16914 8511 16972 8517
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 21174 8440 21180 8492
rect 21232 8480 21238 8492
rect 21453 8483 21511 8489
rect 21453 8480 21465 8483
rect 21232 8452 21465 8480
rect 21232 8440 21238 8452
rect 21453 8449 21465 8452
rect 21499 8449 21511 8483
rect 21453 8443 21511 8449
rect 14001 8415 14059 8421
rect 14001 8412 14013 8415
rect 13556 8384 14013 8412
rect 11517 8375 11575 8381
rect 9582 8304 9588 8356
rect 9640 8344 9646 8356
rect 11054 8344 11060 8356
rect 9640 8316 11060 8344
rect 9640 8304 9646 8316
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 9364 8248 9536 8276
rect 9364 8236 9370 8248
rect 10226 8236 10232 8288
rect 10284 8236 10290 8288
rect 10410 8236 10416 8288
rect 10468 8276 10474 8288
rect 10962 8276 10968 8288
rect 10468 8248 10968 8276
rect 10468 8236 10474 8248
rect 10962 8236 10968 8248
rect 11020 8276 11026 8288
rect 11532 8276 11560 8375
rect 13446 8304 13452 8356
rect 13504 8304 13510 8356
rect 13740 8288 13768 8384
rect 14001 8381 14013 8384
rect 14047 8381 14059 8415
rect 14001 8375 14059 8381
rect 17678 8372 17684 8424
rect 17736 8412 17742 8424
rect 18693 8415 18751 8421
rect 18693 8412 18705 8415
rect 17736 8384 18705 8412
rect 17736 8372 17742 8384
rect 18693 8381 18705 8384
rect 18739 8381 18751 8415
rect 18693 8375 18751 8381
rect 17972 8316 18644 8344
rect 11020 8248 11560 8276
rect 11020 8236 11026 8248
rect 13722 8236 13728 8288
rect 13780 8236 13786 8288
rect 13814 8236 13820 8288
rect 13872 8236 13878 8288
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 15381 8279 15439 8285
rect 15381 8276 15393 8279
rect 15344 8248 15393 8276
rect 15344 8236 15350 8248
rect 15381 8245 15393 8248
rect 15427 8245 15439 8279
rect 15381 8239 15439 8245
rect 15470 8236 15476 8288
rect 15528 8276 15534 8288
rect 16390 8276 16396 8288
rect 15528 8248 16396 8276
rect 15528 8236 15534 8248
rect 16390 8236 16396 8248
rect 16448 8276 16454 8288
rect 17972 8276 18000 8316
rect 18616 8288 18644 8316
rect 16448 8248 18000 8276
rect 16448 8236 16454 8248
rect 18046 8236 18052 8288
rect 18104 8236 18110 8288
rect 18598 8236 18604 8288
rect 18656 8236 18662 8288
rect 1104 8186 22264 8208
rect 1104 8134 3595 8186
rect 3647 8134 3659 8186
rect 3711 8134 3723 8186
rect 3775 8134 3787 8186
rect 3839 8134 3851 8186
rect 3903 8134 8885 8186
rect 8937 8134 8949 8186
rect 9001 8134 9013 8186
rect 9065 8134 9077 8186
rect 9129 8134 9141 8186
rect 9193 8134 14175 8186
rect 14227 8134 14239 8186
rect 14291 8134 14303 8186
rect 14355 8134 14367 8186
rect 14419 8134 14431 8186
rect 14483 8134 19465 8186
rect 19517 8134 19529 8186
rect 19581 8134 19593 8186
rect 19645 8134 19657 8186
rect 19709 8134 19721 8186
rect 19773 8134 22264 8186
rect 1104 8112 22264 8134
rect 6104 8044 7604 8072
rect 6104 8016 6132 8044
rect 6086 7964 6092 8016
rect 6144 7964 6150 8016
rect 7466 8004 7472 8016
rect 7208 7976 7472 8004
rect 6914 7936 6920 7948
rect 5184 7908 6920 7936
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3568 7840 3801 7868
rect 3568 7828 3574 7840
rect 3789 7837 3801 7840
rect 3835 7868 3847 7871
rect 3878 7868 3884 7880
rect 3835 7840 3884 7868
rect 3835 7837 3847 7840
rect 3789 7831 3847 7837
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 4056 7803 4114 7809
rect 4056 7769 4068 7803
rect 4102 7800 4114 7803
rect 4154 7800 4160 7812
rect 4102 7772 4160 7800
rect 4102 7769 4114 7772
rect 4056 7763 4114 7769
rect 4154 7760 4160 7772
rect 4212 7760 4218 7812
rect 5184 7744 5212 7908
rect 6914 7896 6920 7908
rect 6972 7936 6978 7948
rect 7208 7945 7236 7976
rect 7466 7964 7472 7976
rect 7524 7964 7530 8016
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 6972 7908 7205 7936
rect 6972 7896 6978 7908
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5350 7868 5356 7880
rect 5307 7840 5356 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 7098 7828 7104 7880
rect 7156 7828 7162 7880
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7868 7527 7871
rect 7576 7868 7604 8044
rect 7650 8032 7656 8084
rect 7708 8032 7714 8084
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 7800 8044 8033 8072
rect 7800 8032 7806 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 8021 8035 8079 8041
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 9214 8072 9220 8084
rect 8619 8044 9220 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8072 10195 8075
rect 10318 8072 10324 8084
rect 10183 8044 10324 8072
rect 10183 8041 10195 8044
rect 10137 8035 10195 8041
rect 10318 8032 10324 8044
rect 10376 8032 10382 8084
rect 11422 8032 11428 8084
rect 11480 8072 11486 8084
rect 11480 8044 11928 8072
rect 11480 8032 11486 8044
rect 9582 8004 9588 8016
rect 7852 7976 9588 8004
rect 7852 7948 7880 7976
rect 7834 7896 7840 7948
rect 7892 7896 7898 7948
rect 8018 7896 8024 7948
rect 8076 7936 8082 7948
rect 8205 7939 8263 7945
rect 8205 7936 8217 7939
rect 8076 7908 8217 7936
rect 8076 7896 8082 7908
rect 8205 7905 8217 7908
rect 8251 7905 8263 7939
rect 8205 7899 8263 7905
rect 8404 7877 8432 7976
rect 9582 7964 9588 7976
rect 9640 7964 9646 8016
rect 11900 8013 11928 8044
rect 12066 8032 12072 8084
rect 12124 8032 12130 8084
rect 13630 8032 13636 8084
rect 13688 8032 13694 8084
rect 13909 8075 13967 8081
rect 13909 8041 13921 8075
rect 13955 8072 13967 8075
rect 14090 8072 14096 8084
rect 13955 8044 14096 8072
rect 13955 8041 13967 8044
rect 13909 8035 13967 8041
rect 14090 8032 14096 8044
rect 14148 8032 14154 8084
rect 14550 8032 14556 8084
rect 14608 8032 14614 8084
rect 14737 8075 14795 8081
rect 14737 8041 14749 8075
rect 14783 8072 14795 8075
rect 15194 8072 15200 8084
rect 14783 8044 15200 8072
rect 14783 8041 14795 8044
rect 14737 8035 14795 8041
rect 15194 8032 15200 8044
rect 15252 8032 15258 8084
rect 15304 8044 17632 8072
rect 11885 8007 11943 8013
rect 11885 7973 11897 8007
rect 11931 8004 11943 8007
rect 13648 8004 13676 8032
rect 11931 7976 13676 8004
rect 11931 7973 11943 7976
rect 11885 7967 11943 7973
rect 13814 7964 13820 8016
rect 13872 7964 13878 8016
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10318 7936 10324 7948
rect 10008 7908 10324 7936
rect 10008 7896 10014 7908
rect 10318 7896 10324 7908
rect 10376 7936 10382 7948
rect 13832 7936 13860 7964
rect 14568 7936 14596 8032
rect 10376 7908 10640 7936
rect 10376 7896 10382 7908
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 7515 7840 7757 7868
rect 7515 7837 7527 7840
rect 7469 7831 7527 7837
rect 7745 7837 7757 7840
rect 7791 7837 7803 7871
rect 8389 7871 8447 7877
rect 7745 7831 7803 7837
rect 7852 7840 8340 7868
rect 6822 7760 6828 7812
rect 6880 7800 6886 7812
rect 7392 7800 7420 7831
rect 7852 7800 7880 7840
rect 6880 7772 7880 7800
rect 6880 7760 6886 7772
rect 8018 7760 8024 7812
rect 8076 7809 8082 7812
rect 8076 7803 8089 7809
rect 8077 7800 8089 7803
rect 8312 7800 8340 7840
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7868 9919 7871
rect 10042 7868 10048 7880
rect 9907 7840 10048 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10134 7828 10140 7880
rect 10192 7828 10198 7880
rect 10226 7828 10232 7880
rect 10284 7828 10290 7880
rect 10410 7828 10416 7880
rect 10468 7868 10474 7880
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 10468 7840 10517 7868
rect 10468 7828 10474 7840
rect 10505 7837 10517 7840
rect 10551 7837 10563 7871
rect 10612 7868 10640 7908
rect 12820 7908 13860 7936
rect 14292 7908 14596 7936
rect 12342 7868 12348 7880
rect 10612 7840 12348 7868
rect 10505 7831 10563 7837
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 12434 7828 12440 7880
rect 12492 7828 12498 7880
rect 12526 7828 12532 7880
rect 12584 7828 12590 7880
rect 12618 7828 12624 7880
rect 12676 7828 12682 7880
rect 12820 7877 12848 7908
rect 14292 7877 14320 7908
rect 15304 7877 15332 8044
rect 17604 8004 17632 8044
rect 17678 8032 17684 8084
rect 17736 8032 17742 8084
rect 18966 8004 18972 8016
rect 17604 7976 18972 8004
rect 18966 7964 18972 7976
rect 19024 7964 19030 8016
rect 15378 7896 15384 7948
rect 15436 7936 15442 7948
rect 16301 7939 16359 7945
rect 16301 7936 16313 7939
rect 15436 7908 16313 7936
rect 15436 7896 15442 7908
rect 16301 7905 16313 7908
rect 16347 7905 16359 7939
rect 16301 7899 16359 7905
rect 18046 7896 18052 7948
rect 18104 7896 18110 7948
rect 21085 7939 21143 7945
rect 21085 7905 21097 7939
rect 21131 7936 21143 7939
rect 21545 7939 21603 7945
rect 21545 7936 21557 7939
rect 21131 7908 21557 7936
rect 21131 7905 21143 7908
rect 21085 7899 21143 7905
rect 21545 7905 21557 7908
rect 21591 7905 21603 7939
rect 21545 7899 21603 7905
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7868 13783 7871
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13771 7840 14105 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 14599 7840 15117 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 10244 7800 10272 7828
rect 10750 7803 10808 7809
rect 10750 7800 10762 7803
rect 8077 7772 8248 7800
rect 8312 7772 10088 7800
rect 10244 7772 10762 7800
rect 8077 7769 8089 7772
rect 8076 7763 8089 7769
rect 8076 7760 8082 7763
rect 5166 7692 5172 7744
rect 5224 7692 5230 7744
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 6549 7735 6607 7741
rect 6549 7732 6561 7735
rect 5592 7704 6561 7732
rect 5592 7692 5598 7704
rect 6549 7701 6561 7704
rect 6595 7701 6607 7735
rect 6549 7695 6607 7701
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7837 7735 7895 7741
rect 7837 7732 7849 7735
rect 6972 7704 7849 7732
rect 6972 7692 6978 7704
rect 7837 7701 7849 7704
rect 7883 7701 7895 7735
rect 8220 7732 8248 7772
rect 8754 7732 8760 7744
rect 8220 7704 8760 7732
rect 7837 7695 7895 7701
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 9953 7735 10011 7741
rect 9953 7732 9965 7735
rect 9916 7704 9965 7732
rect 9916 7692 9922 7704
rect 9953 7701 9965 7704
rect 9999 7701 10011 7735
rect 10060 7732 10088 7772
rect 10750 7769 10762 7772
rect 10796 7769 10808 7803
rect 10750 7763 10808 7769
rect 11974 7760 11980 7812
rect 12032 7800 12038 7812
rect 12820 7800 12848 7831
rect 12032 7772 12848 7800
rect 14476 7800 14504 7831
rect 15470 7828 15476 7880
rect 15528 7828 15534 7880
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7868 16083 7871
rect 16071 7840 16712 7868
rect 16071 7837 16083 7840
rect 16025 7831 16083 7837
rect 16684 7812 16712 7840
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19429 7871 19487 7877
rect 19429 7868 19441 7871
rect 19392 7840 19441 7868
rect 19392 7828 19398 7840
rect 19429 7837 19441 7840
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 20533 7871 20591 7877
rect 20533 7837 20545 7871
rect 20579 7868 20591 7871
rect 20622 7868 20628 7880
rect 20579 7840 20628 7868
rect 20579 7837 20591 7840
rect 20533 7831 20591 7837
rect 16546 7803 16604 7809
rect 16546 7800 16558 7803
rect 14476 7772 14596 7800
rect 12032 7760 12038 7772
rect 11992 7732 12020 7760
rect 14568 7744 14596 7772
rect 16224 7772 16558 7800
rect 10060 7704 12020 7732
rect 9953 7695 10011 7701
rect 14550 7692 14556 7744
rect 14608 7692 14614 7744
rect 16224 7741 16252 7772
rect 16546 7769 16558 7772
rect 16592 7769 16604 7803
rect 16546 7763 16604 7769
rect 16666 7760 16672 7812
rect 16724 7760 16730 7812
rect 20180 7800 20208 7831
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 20772 7840 21373 7868
rect 20772 7828 20778 7840
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 21818 7828 21824 7880
rect 21876 7828 21882 7880
rect 21177 7803 21235 7809
rect 21177 7800 21189 7803
rect 20180 7772 21189 7800
rect 21177 7769 21189 7772
rect 21223 7769 21235 7803
rect 21177 7763 21235 7769
rect 16209 7735 16267 7741
rect 16209 7701 16221 7735
rect 16255 7701 16267 7735
rect 16209 7695 16267 7701
rect 18414 7692 18420 7744
rect 18472 7732 18478 7744
rect 18693 7735 18751 7741
rect 18693 7732 18705 7735
rect 18472 7704 18705 7732
rect 18472 7692 18478 7704
rect 18693 7701 18705 7704
rect 18739 7701 18751 7735
rect 18693 7695 18751 7701
rect 19242 7692 19248 7744
rect 19300 7692 19306 7744
rect 20349 7735 20407 7741
rect 20349 7701 20361 7735
rect 20395 7732 20407 7735
rect 20806 7732 20812 7744
rect 20395 7704 20812 7732
rect 20395 7701 20407 7704
rect 20349 7695 20407 7701
rect 20806 7692 20812 7704
rect 20864 7692 20870 7744
rect 21542 7692 21548 7744
rect 21600 7732 21606 7744
rect 21637 7735 21695 7741
rect 21637 7732 21649 7735
rect 21600 7704 21649 7732
rect 21600 7692 21606 7704
rect 21637 7701 21649 7704
rect 21683 7701 21695 7735
rect 21637 7695 21695 7701
rect 1104 7642 22264 7664
rect 1104 7590 4255 7642
rect 4307 7590 4319 7642
rect 4371 7590 4383 7642
rect 4435 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 9545 7642
rect 9597 7590 9609 7642
rect 9661 7590 9673 7642
rect 9725 7590 9737 7642
rect 9789 7590 9801 7642
rect 9853 7590 14835 7642
rect 14887 7590 14899 7642
rect 14951 7590 14963 7642
rect 15015 7590 15027 7642
rect 15079 7590 15091 7642
rect 15143 7590 20125 7642
rect 20177 7590 20189 7642
rect 20241 7590 20253 7642
rect 20305 7590 20317 7642
rect 20369 7590 20381 7642
rect 20433 7590 22264 7642
rect 1104 7568 22264 7590
rect 5074 7488 5080 7540
rect 5132 7528 5138 7540
rect 5563 7531 5621 7537
rect 5132 7500 5396 7528
rect 5132 7488 5138 7500
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 5258 7460 5264 7472
rect 4387 7432 5264 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 5258 7420 5264 7432
rect 5316 7420 5322 7472
rect 5368 7469 5396 7500
rect 5563 7497 5575 7531
rect 5609 7528 5621 7531
rect 6086 7528 6092 7540
rect 5609 7500 6092 7528
rect 5609 7497 5621 7500
rect 5563 7491 5621 7497
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 6457 7531 6515 7537
rect 6457 7497 6469 7531
rect 6503 7528 6515 7531
rect 7006 7528 7012 7540
rect 6503 7500 7012 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 11517 7531 11575 7537
rect 7156 7500 7328 7528
rect 7156 7488 7162 7500
rect 5353 7463 5411 7469
rect 5353 7429 5365 7463
rect 5399 7429 5411 7463
rect 5353 7423 5411 7429
rect 5166 7352 5172 7404
rect 5224 7352 5230 7404
rect 3053 7191 3111 7197
rect 3053 7157 3065 7191
rect 3099 7188 3111 7191
rect 3970 7188 3976 7200
rect 3099 7160 3976 7188
rect 3099 7157 3111 7160
rect 3053 7151 3111 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 5184 7188 5212 7352
rect 5368 7324 5396 7423
rect 6104 7392 6132 7488
rect 6822 7420 6828 7472
rect 6880 7420 6886 7472
rect 7300 7460 7328 7500
rect 11517 7497 11529 7531
rect 11563 7528 11575 7531
rect 11698 7528 11704 7540
rect 11563 7500 11704 7528
rect 11563 7497 11575 7500
rect 11517 7491 11575 7497
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 11974 7488 11980 7540
rect 12032 7488 12038 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 13909 7531 13967 7537
rect 13909 7528 13921 7531
rect 12492 7500 13921 7528
rect 12492 7488 12498 7500
rect 13909 7497 13921 7500
rect 13955 7497 13967 7531
rect 19521 7531 19579 7537
rect 19521 7528 19533 7531
rect 13909 7491 13967 7497
rect 19352 7500 19533 7528
rect 8021 7463 8079 7469
rect 8021 7460 8033 7463
rect 7300 7432 8033 7460
rect 6641 7395 6699 7401
rect 6641 7392 6653 7395
rect 6104 7364 6653 7392
rect 6641 7361 6653 7364
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 6840 7392 6868 7420
rect 6779 7364 6868 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 6914 7352 6920 7404
rect 6972 7352 6978 7404
rect 7019 7385 7077 7391
rect 6932 7324 6960 7352
rect 7019 7351 7031 7385
rect 7065 7351 7077 7385
rect 7282 7352 7288 7404
rect 7340 7352 7346 7404
rect 7374 7352 7380 7404
rect 7432 7352 7438 7404
rect 7466 7352 7472 7404
rect 7524 7352 7530 7404
rect 7668 7401 7696 7432
rect 8021 7429 8033 7432
rect 8067 7429 8079 7463
rect 8021 7423 8079 7429
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 8386 7392 8392 7404
rect 8159 7364 8392 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7392 11943 7395
rect 11992 7392 12020 7488
rect 14550 7460 14556 7472
rect 14016 7432 14556 7460
rect 11931 7364 12020 7392
rect 13817 7395 13875 7401
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 13817 7361 13829 7395
rect 13863 7392 13875 7395
rect 13906 7392 13912 7404
rect 13863 7364 13912 7392
rect 13863 7361 13875 7364
rect 13817 7355 13875 7361
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 14016 7401 14044 7432
rect 14550 7420 14556 7432
rect 14608 7460 14614 7472
rect 19352 7460 19380 7500
rect 19521 7497 19533 7500
rect 19567 7497 19579 7531
rect 19521 7491 19579 7497
rect 20257 7531 20315 7537
rect 20257 7497 20269 7531
rect 20303 7528 20315 7531
rect 20622 7528 20628 7540
rect 20303 7500 20628 7528
rect 20303 7497 20315 7500
rect 20257 7491 20315 7497
rect 19978 7460 19984 7472
rect 14608 7432 19380 7460
rect 19812 7432 19984 7460
rect 14608 7420 14614 7432
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14642 7392 14648 7404
rect 14507 7364 14648 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 17773 7395 17831 7401
rect 17773 7361 17785 7395
rect 17819 7361 17831 7395
rect 17773 7355 17831 7361
rect 17957 7395 18015 7401
rect 17957 7361 17969 7395
rect 18003 7392 18015 7395
rect 18233 7395 18291 7401
rect 18003 7364 18184 7392
rect 18003 7361 18015 7364
rect 17957 7355 18015 7361
rect 7019 7345 7077 7351
rect 5368 7296 6960 7324
rect 5537 7191 5595 7197
rect 5537 7188 5549 7191
rect 5184 7160 5549 7188
rect 5537 7157 5549 7160
rect 5583 7157 5595 7191
rect 5537 7151 5595 7157
rect 5718 7148 5724 7200
rect 5776 7148 5782 7200
rect 7034 7188 7062 7345
rect 8294 7324 8300 7336
rect 7116 7296 8300 7324
rect 7116 7265 7144 7296
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12066 7324 12072 7336
rect 12023 7296 12072 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 12066 7284 12072 7296
rect 12124 7284 12130 7336
rect 14737 7327 14795 7333
rect 14737 7293 14749 7327
rect 14783 7324 14795 7327
rect 15286 7324 15292 7336
rect 14783 7296 15292 7324
rect 14783 7293 14795 7296
rect 14737 7287 14795 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 17494 7284 17500 7336
rect 17552 7284 17558 7336
rect 17788 7324 17816 7355
rect 18046 7324 18052 7336
rect 17788 7296 18052 7324
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 7101 7259 7159 7265
rect 7101 7225 7113 7259
rect 7147 7225 7159 7259
rect 7101 7219 7159 7225
rect 10318 7188 10324 7200
rect 7034 7160 10324 7188
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 14093 7191 14151 7197
rect 14093 7188 14105 7191
rect 12676 7160 14105 7188
rect 12676 7148 12682 7160
rect 14093 7157 14105 7160
rect 14139 7157 14151 7191
rect 14093 7151 14151 7157
rect 16853 7191 16911 7197
rect 16853 7157 16865 7191
rect 16899 7188 16911 7191
rect 16942 7188 16948 7200
rect 16899 7160 16948 7188
rect 16899 7157 16911 7160
rect 16853 7151 16911 7157
rect 16942 7148 16948 7160
rect 17000 7148 17006 7200
rect 18156 7188 18184 7364
rect 18233 7361 18245 7395
rect 18279 7392 18291 7395
rect 18785 7395 18843 7401
rect 18785 7392 18797 7395
rect 18279 7364 18797 7392
rect 18279 7361 18291 7364
rect 18233 7355 18291 7361
rect 18785 7361 18797 7364
rect 18831 7392 18843 7395
rect 19242 7392 19248 7404
rect 18831 7364 19248 7392
rect 18831 7361 18843 7364
rect 18785 7355 18843 7361
rect 19242 7352 19248 7364
rect 19300 7352 19306 7404
rect 19812 7401 19840 7432
rect 19978 7420 19984 7432
rect 20036 7460 20042 7472
rect 20272 7460 20300 7491
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 20036 7432 20300 7460
rect 20036 7420 20042 7432
rect 20530 7420 20536 7472
rect 20588 7460 20594 7472
rect 20588 7432 21680 7460
rect 20588 7420 20594 7432
rect 19797 7395 19855 7401
rect 19797 7361 19809 7395
rect 19843 7361 19855 7395
rect 19797 7355 19855 7361
rect 20073 7395 20131 7401
rect 20073 7361 20085 7395
rect 20119 7392 20131 7395
rect 20162 7392 20168 7404
rect 20119 7364 20168 7392
rect 20119 7361 20131 7364
rect 20073 7355 20131 7361
rect 20162 7352 20168 7364
rect 20220 7392 20226 7404
rect 20622 7392 20628 7404
rect 20220 7364 20628 7392
rect 20220 7352 20226 7364
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 21381 7395 21439 7401
rect 21381 7361 21393 7395
rect 21427 7392 21439 7395
rect 21542 7392 21548 7404
rect 21427 7364 21548 7392
rect 21427 7361 21439 7364
rect 21381 7355 21439 7361
rect 21542 7352 21548 7364
rect 21600 7352 21606 7404
rect 21652 7401 21680 7432
rect 21637 7395 21695 7401
rect 21637 7361 21649 7395
rect 21683 7361 21695 7395
rect 21637 7355 21695 7361
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 18463 7296 18521 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 18509 7293 18521 7296
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 19886 7284 19892 7336
rect 19944 7284 19950 7336
rect 19613 7259 19671 7265
rect 19613 7256 19625 7259
rect 19076 7228 19625 7256
rect 19076 7188 19104 7228
rect 19613 7225 19625 7228
rect 19659 7225 19671 7259
rect 19613 7219 19671 7225
rect 18156 7160 19104 7188
rect 20073 7191 20131 7197
rect 20073 7157 20085 7191
rect 20119 7188 20131 7191
rect 20438 7188 20444 7200
rect 20119 7160 20444 7188
rect 20119 7157 20131 7160
rect 20073 7151 20131 7157
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 1104 7098 22264 7120
rect 1104 7046 3595 7098
rect 3647 7046 3659 7098
rect 3711 7046 3723 7098
rect 3775 7046 3787 7098
rect 3839 7046 3851 7098
rect 3903 7046 8885 7098
rect 8937 7046 8949 7098
rect 9001 7046 9013 7098
rect 9065 7046 9077 7098
rect 9129 7046 9141 7098
rect 9193 7046 14175 7098
rect 14227 7046 14239 7098
rect 14291 7046 14303 7098
rect 14355 7046 14367 7098
rect 14419 7046 14431 7098
rect 14483 7046 19465 7098
rect 19517 7046 19529 7098
rect 19581 7046 19593 7098
rect 19645 7046 19657 7098
rect 19709 7046 19721 7098
rect 19773 7046 22264 7098
rect 1104 7024 22264 7046
rect 8018 6944 8024 6996
rect 8076 6984 8082 6996
rect 8076 6956 10824 6984
rect 8076 6944 8082 6956
rect 9585 6919 9643 6925
rect 9585 6885 9597 6919
rect 9631 6916 9643 6919
rect 9631 6888 10088 6916
rect 9631 6885 9643 6888
rect 9585 6879 9643 6885
rect 4801 6851 4859 6857
rect 4801 6817 4813 6851
rect 4847 6848 4859 6851
rect 4847 6820 5304 6848
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 5276 6789 5304 6820
rect 7190 6808 7196 6860
rect 7248 6848 7254 6860
rect 8478 6848 8484 6860
rect 7248 6820 8484 6848
rect 7248 6808 7254 6820
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 9858 6848 9864 6860
rect 9048 6820 9864 6848
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4120 6752 5089 6780
rect 4120 6740 4126 6752
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6780 5319 6783
rect 7282 6780 7288 6792
rect 5307 6752 7288 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5092 6712 5120 6743
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 8018 6740 8024 6792
rect 8076 6740 8082 6792
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6780 8355 6783
rect 8570 6780 8576 6792
rect 8343 6752 8576 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 9048 6789 9076 6820
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 10060 6857 10088 6888
rect 10045 6851 10103 6857
rect 10045 6817 10057 6851
rect 10091 6817 10103 6851
rect 10708 6851 10766 6857
rect 10708 6848 10720 6851
rect 10045 6811 10103 6817
rect 10244 6820 10720 6848
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 8680 6752 9045 6780
rect 5718 6712 5724 6724
rect 5092 6684 5724 6712
rect 5718 6672 5724 6684
rect 5776 6712 5782 6724
rect 6454 6712 6460 6724
rect 5776 6684 6460 6712
rect 5776 6672 5782 6684
rect 6454 6672 6460 6684
rect 6512 6672 6518 6724
rect 8202 6672 8208 6724
rect 8260 6672 8266 6724
rect 8680 6656 8708 6752
rect 9033 6749 9045 6752
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 9214 6740 9220 6792
rect 9272 6740 9278 6792
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 9456 6752 9505 6780
rect 9456 6740 9462 6752
rect 9493 6749 9505 6752
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6749 10011 6783
rect 9953 6743 10011 6749
rect 9858 6672 9864 6724
rect 9916 6672 9922 6724
rect 4154 6604 4160 6656
rect 4212 6604 4218 6656
rect 4890 6604 4896 6656
rect 4948 6604 4954 6656
rect 8119 6647 8177 6653
rect 8119 6613 8131 6647
rect 8165 6644 8177 6647
rect 8386 6644 8392 6656
rect 8165 6616 8392 6644
rect 8165 6613 8177 6616
rect 8119 6607 8177 6613
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 8662 6604 8668 6656
rect 8720 6604 8726 6656
rect 9968 6644 9996 6743
rect 10060 6712 10088 6811
rect 10244 6789 10272 6820
rect 10708 6817 10720 6820
rect 10754 6817 10766 6851
rect 10708 6811 10766 6817
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 10410 6740 10416 6792
rect 10468 6740 10474 6792
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 10520 6712 10548 6743
rect 10796 6721 10824 6956
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 13449 6987 13507 6993
rect 13449 6984 13461 6987
rect 12584 6956 13461 6984
rect 12584 6944 12590 6956
rect 13449 6953 13461 6956
rect 13495 6953 13507 6987
rect 13449 6947 13507 6953
rect 16666 6944 16672 6996
rect 16724 6944 16730 6996
rect 17586 6944 17592 6996
rect 17644 6984 17650 6996
rect 17954 6984 17960 6996
rect 17644 6956 17960 6984
rect 17644 6944 17650 6956
rect 17954 6944 17960 6956
rect 18012 6944 18018 6996
rect 18046 6944 18052 6996
rect 18104 6984 18110 6996
rect 18233 6987 18291 6993
rect 18233 6984 18245 6987
rect 18104 6956 18245 6984
rect 18104 6944 18110 6956
rect 18233 6953 18245 6956
rect 18279 6953 18291 6987
rect 18233 6947 18291 6953
rect 19245 6987 19303 6993
rect 19245 6953 19257 6987
rect 19291 6984 19303 6987
rect 19334 6984 19340 6996
rect 19291 6956 19340 6984
rect 19291 6953 19303 6956
rect 19245 6947 19303 6953
rect 19334 6944 19340 6956
rect 19392 6944 19398 6996
rect 19429 6987 19487 6993
rect 19429 6953 19441 6987
rect 19475 6953 19487 6987
rect 19429 6947 19487 6953
rect 13633 6919 13691 6925
rect 13633 6885 13645 6919
rect 13679 6885 13691 6919
rect 13633 6879 13691 6885
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11204 6820 11989 6848
rect 11204 6808 11210 6820
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 13648 6848 13676 6879
rect 17678 6876 17684 6928
rect 17736 6876 17742 6928
rect 17788 6888 18000 6916
rect 13906 6848 13912 6860
rect 13648 6820 13912 6848
rect 11977 6811 12035 6817
rect 13906 6808 13912 6820
rect 13964 6848 13970 6860
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 13964 6820 14657 6848
rect 13964 6808 13970 6820
rect 14645 6817 14657 6820
rect 14691 6817 14703 6851
rect 16114 6848 16120 6860
rect 14645 6811 14703 6817
rect 15304 6820 16120 6848
rect 11701 6783 11759 6789
rect 11701 6749 11713 6783
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 10060 6684 10548 6712
rect 10781 6715 10839 6721
rect 10781 6681 10793 6715
rect 10827 6681 10839 6715
rect 11716 6712 11744 6743
rect 11882 6740 11888 6792
rect 11940 6740 11946 6792
rect 12066 6740 12072 6792
rect 12124 6740 12130 6792
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6780 14519 6783
rect 14550 6780 14556 6792
rect 14507 6752 14556 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 15304 6789 15332 6820
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 17129 6851 17187 6857
rect 17129 6817 17141 6851
rect 17175 6848 17187 6851
rect 17788 6848 17816 6888
rect 17175 6820 17816 6848
rect 17175 6817 17187 6820
rect 17129 6811 17187 6817
rect 17862 6808 17868 6860
rect 17920 6808 17926 6860
rect 17972 6848 18000 6888
rect 19444 6848 19472 6947
rect 19886 6944 19892 6996
rect 19944 6944 19950 6996
rect 17972 6820 19472 6848
rect 20530 6808 20536 6860
rect 20588 6808 20594 6860
rect 15105 6783 15163 6789
rect 15105 6780 15117 6783
rect 14660 6752 15117 6780
rect 12084 6712 12112 6740
rect 11716 6684 12112 6712
rect 13909 6715 13967 6721
rect 10781 6675 10839 6681
rect 13909 6681 13921 6715
rect 13955 6712 13967 6715
rect 14660 6712 14688 6752
rect 15105 6749 15117 6752
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 16301 6783 16359 6789
rect 16301 6780 16313 6783
rect 15896 6752 16313 6780
rect 15896 6740 15902 6752
rect 16301 6749 16313 6752
rect 16347 6749 16359 6783
rect 16301 6743 16359 6749
rect 16850 6740 16856 6792
rect 16908 6740 16914 6792
rect 16942 6740 16948 6792
rect 17000 6740 17006 6792
rect 17313 6783 17371 6789
rect 17313 6749 17325 6783
rect 17359 6780 17371 6783
rect 17494 6780 17500 6792
rect 17359 6752 17500 6780
rect 17359 6749 17371 6752
rect 17313 6743 17371 6749
rect 17494 6740 17500 6752
rect 17552 6780 17558 6792
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 17552 6752 17816 6780
rect 17552 6740 17558 6752
rect 17586 6712 17592 6724
rect 13955 6684 14688 6712
rect 13955 6681 13967 6684
rect 13909 6675 13967 6681
rect 14660 6656 14688 6684
rect 17512 6684 17592 6712
rect 10042 6644 10048 6656
rect 9968 6616 10048 6644
rect 10042 6604 10048 6616
rect 10100 6644 10106 6656
rect 10597 6647 10655 6653
rect 10597 6644 10609 6647
rect 10100 6616 10609 6644
rect 10100 6604 10106 6616
rect 10597 6613 10609 6616
rect 10643 6613 10655 6647
rect 10597 6607 10655 6613
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 14553 6647 14611 6653
rect 14553 6613 14565 6647
rect 14599 6644 14611 6647
rect 14642 6644 14648 6656
rect 14599 6616 14648 6644
rect 14599 6613 14611 6616
rect 14553 6607 14611 6613
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 15470 6604 15476 6656
rect 15528 6604 15534 6656
rect 16485 6647 16543 6653
rect 16485 6613 16497 6647
rect 16531 6644 16543 6647
rect 16850 6644 16856 6656
rect 16531 6616 16856 6644
rect 16531 6613 16543 6616
rect 16485 6607 16543 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 17402 6604 17408 6656
rect 17460 6604 17466 6656
rect 17512 6653 17540 6684
rect 17586 6672 17592 6684
rect 17644 6672 17650 6724
rect 17678 6672 17684 6724
rect 17736 6672 17742 6724
rect 17788 6721 17816 6752
rect 17972 6752 18061 6780
rect 17773 6715 17831 6721
rect 17773 6681 17785 6715
rect 17819 6712 17831 6715
rect 17862 6712 17868 6724
rect 17819 6684 17868 6712
rect 17819 6681 17831 6684
rect 17773 6675 17831 6681
rect 17862 6672 17868 6684
rect 17920 6672 17926 6724
rect 17497 6647 17555 6653
rect 17497 6613 17509 6647
rect 17543 6613 17555 6647
rect 17696 6644 17724 6672
rect 17972 6644 18000 6752
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 18414 6740 18420 6792
rect 18472 6740 18478 6792
rect 20806 6789 20812 6792
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6749 18567 6783
rect 18509 6743 18567 6749
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6780 18751 6783
rect 18969 6783 19027 6789
rect 18969 6780 18981 6783
rect 18739 6752 18981 6780
rect 18739 6749 18751 6752
rect 18693 6743 18751 6749
rect 18969 6749 18981 6752
rect 19015 6749 19027 6783
rect 20800 6780 20812 6789
rect 18969 6743 19027 6749
rect 19628 6752 20484 6780
rect 20767 6752 20812 6780
rect 18524 6712 18552 6743
rect 19628 6721 19656 6752
rect 18064 6684 18552 6712
rect 19613 6715 19671 6721
rect 18064 6656 18092 6684
rect 19613 6681 19625 6715
rect 19659 6681 19671 6715
rect 19613 6675 19671 6681
rect 19978 6672 19984 6724
rect 20036 6712 20042 6724
rect 20073 6715 20131 6721
rect 20073 6712 20085 6715
rect 20036 6684 20085 6712
rect 20036 6672 20042 6684
rect 20073 6681 20085 6684
rect 20119 6681 20131 6715
rect 20073 6675 20131 6681
rect 20456 6656 20484 6752
rect 20800 6743 20812 6752
rect 20806 6740 20812 6743
rect 20864 6740 20870 6792
rect 17696 6616 18000 6644
rect 17497 6607 17555 6613
rect 18046 6604 18052 6656
rect 18104 6604 18110 6656
rect 18782 6604 18788 6656
rect 18840 6604 18846 6656
rect 19413 6647 19471 6653
rect 19413 6613 19425 6647
rect 19459 6644 19471 6647
rect 19705 6647 19763 6653
rect 19705 6644 19717 6647
rect 19459 6616 19717 6644
rect 19459 6613 19471 6616
rect 19413 6607 19471 6613
rect 19705 6613 19717 6616
rect 19751 6613 19763 6647
rect 19705 6607 19763 6613
rect 19873 6647 19931 6653
rect 19873 6613 19885 6647
rect 19919 6644 19931 6647
rect 20162 6644 20168 6656
rect 19919 6616 20168 6644
rect 19919 6613 19931 6616
rect 19873 6607 19931 6613
rect 20162 6604 20168 6616
rect 20220 6604 20226 6656
rect 20438 6604 20444 6656
rect 20496 6644 20502 6656
rect 21913 6647 21971 6653
rect 21913 6644 21925 6647
rect 20496 6616 21925 6644
rect 20496 6604 20502 6616
rect 21913 6613 21925 6616
rect 21959 6613 21971 6647
rect 21913 6607 21971 6613
rect 1104 6554 22264 6576
rect 1104 6502 4255 6554
rect 4307 6502 4319 6554
rect 4371 6502 4383 6554
rect 4435 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 9545 6554
rect 9597 6502 9609 6554
rect 9661 6502 9673 6554
rect 9725 6502 9737 6554
rect 9789 6502 9801 6554
rect 9853 6502 14835 6554
rect 14887 6502 14899 6554
rect 14951 6502 14963 6554
rect 15015 6502 15027 6554
rect 15079 6502 15091 6554
rect 15143 6502 20125 6554
rect 20177 6502 20189 6554
rect 20241 6502 20253 6554
rect 20305 6502 20317 6554
rect 20369 6502 20381 6554
rect 20433 6502 22264 6554
rect 1104 6480 22264 6502
rect 4062 6400 4068 6452
rect 4120 6400 4126 6452
rect 4154 6400 4160 6452
rect 4212 6400 4218 6452
rect 7190 6440 7196 6452
rect 4908 6412 5856 6440
rect 4080 6372 4108 6400
rect 3988 6344 4108 6372
rect 3988 6313 4016 6344
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6273 4031 6307
rect 3973 6267 4031 6273
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6304 4123 6307
rect 4172 6304 4200 6400
rect 4908 6384 4936 6412
rect 4890 6332 4896 6384
rect 4948 6332 4954 6384
rect 5292 6375 5350 6381
rect 5292 6341 5304 6375
rect 5338 6372 5350 6375
rect 5721 6375 5779 6381
rect 5721 6372 5733 6375
rect 5338 6344 5733 6372
rect 5338 6341 5350 6344
rect 5292 6335 5350 6341
rect 5721 6341 5733 6344
rect 5767 6341 5779 6375
rect 5721 6335 5779 6341
rect 5828 6313 5856 6412
rect 6564 6412 7196 6440
rect 6564 6313 6592 6412
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 7282 6400 7288 6452
rect 7340 6400 7346 6452
rect 8386 6400 8392 6452
rect 8444 6400 8450 6452
rect 8570 6400 8576 6452
rect 8628 6400 8634 6452
rect 9214 6400 9220 6452
rect 9272 6400 9278 6452
rect 9861 6443 9919 6449
rect 9861 6409 9873 6443
rect 9907 6440 9919 6443
rect 10042 6440 10048 6452
rect 9907 6412 10048 6440
rect 9907 6409 9919 6412
rect 9861 6403 9919 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10410 6400 10416 6452
rect 10468 6400 10474 6452
rect 11514 6400 11520 6452
rect 11572 6440 11578 6452
rect 11701 6443 11759 6449
rect 11701 6440 11713 6443
rect 11572 6412 11713 6440
rect 11572 6400 11578 6412
rect 11701 6409 11713 6412
rect 11747 6409 11759 6443
rect 11701 6403 11759 6409
rect 11882 6400 11888 6452
rect 11940 6440 11946 6452
rect 13173 6443 13231 6449
rect 13173 6440 13185 6443
rect 11940 6412 13185 6440
rect 11940 6400 11946 6412
rect 7300 6372 7328 6400
rect 6748 6344 7328 6372
rect 6748 6313 6776 6344
rect 8018 6332 8024 6384
rect 8076 6372 8082 6384
rect 8205 6375 8263 6381
rect 8205 6372 8217 6375
rect 8076 6344 8217 6372
rect 8076 6332 8082 6344
rect 8205 6341 8217 6344
rect 8251 6341 8263 6375
rect 8205 6335 8263 6341
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 4111 6276 4200 6304
rect 4540 6276 5641 6304
rect 4111 6273 4123 6276
rect 4065 6267 4123 6273
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 3789 6239 3847 6245
rect 3789 6236 3801 6239
rect 3292 6208 3801 6236
rect 3292 6196 3298 6208
rect 3789 6205 3801 6208
rect 3835 6205 3847 6239
rect 3789 6199 3847 6205
rect 3881 6171 3939 6177
rect 3881 6137 3893 6171
rect 3927 6168 3939 6171
rect 4540 6168 4568 6276
rect 5629 6273 5641 6276
rect 5675 6273 5687 6307
rect 5629 6267 5687 6273
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6304 6883 6307
rect 6871 6276 7052 6304
rect 6871 6273 6883 6276
rect 6825 6267 6883 6273
rect 5534 6196 5540 6248
rect 5592 6196 5598 6248
rect 3927 6140 4568 6168
rect 3927 6137 3939 6140
rect 3881 6131 3939 6137
rect 4157 6103 4215 6109
rect 4157 6069 4169 6103
rect 4203 6100 4215 6103
rect 6748 6100 6776 6267
rect 6914 6196 6920 6248
rect 6972 6196 6978 6248
rect 7024 6236 7052 6276
rect 7098 6264 7104 6316
rect 7156 6264 7162 6316
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 8404 6313 8432 6400
rect 8588 6313 8616 6400
rect 10220 6375 10278 6381
rect 8680 6344 9904 6372
rect 8680 6313 8708 6344
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 7616 6276 7757 6304
rect 7616 6264 7622 6276
rect 7745 6273 7757 6276
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 7374 6236 7380 6248
rect 7024 6208 7380 6236
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7834 6196 7840 6248
rect 7892 6196 7898 6248
rect 8202 6236 8208 6248
rect 8128 6208 8208 6236
rect 4203 6072 6776 6100
rect 7285 6103 7343 6109
rect 4203 6069 4215 6072
rect 4157 6063 4215 6069
rect 7285 6069 7297 6103
rect 7331 6100 7343 6103
rect 7374 6100 7380 6112
rect 7331 6072 7380 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 7852 6100 7880 6196
rect 8128 6177 8156 6208
rect 8202 6196 8208 6208
rect 8260 6236 8266 6248
rect 8680 6236 8708 6267
rect 8754 6264 8760 6316
rect 8812 6304 8818 6316
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8812 6276 8861 6304
rect 8812 6264 8818 6276
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6304 9091 6307
rect 9079 6276 9260 6304
rect 9079 6273 9091 6276
rect 9033 6267 9091 6273
rect 9232 6248 9260 6276
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 9364 6276 9505 6304
rect 9364 6264 9370 6276
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 9876 6248 9904 6344
rect 10220 6341 10232 6375
rect 10266 6372 10278 6375
rect 10428 6372 10456 6400
rect 12360 6381 12388 6412
rect 13173 6409 13185 6412
rect 13219 6409 13231 6443
rect 13173 6403 13231 6409
rect 13906 6400 13912 6452
rect 13964 6400 13970 6452
rect 14090 6400 14096 6452
rect 14148 6400 14154 6452
rect 15381 6443 15439 6449
rect 15381 6409 15393 6443
rect 15427 6409 15439 6443
rect 15381 6403 15439 6409
rect 10266 6344 10456 6372
rect 12345 6375 12403 6381
rect 10266 6341 10278 6344
rect 10220 6335 10278 6341
rect 12345 6341 12357 6375
rect 12391 6372 12403 6375
rect 12391 6344 12425 6372
rect 12391 6341 12403 6344
rect 12345 6335 12403 6341
rect 12618 6332 12624 6384
rect 12676 6372 12682 6384
rect 13262 6372 13268 6384
rect 12676 6344 13268 6372
rect 12676 6332 12682 6344
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 13633 6375 13691 6381
rect 13633 6341 13645 6375
rect 13679 6372 13691 6375
rect 14108 6372 14136 6400
rect 13679 6344 14136 6372
rect 15044 6375 15102 6381
rect 13679 6341 13691 6344
rect 13633 6335 13691 6341
rect 15044 6341 15056 6375
rect 15090 6372 15102 6375
rect 15396 6372 15424 6403
rect 15470 6400 15476 6452
rect 15528 6400 15534 6452
rect 17402 6440 17408 6452
rect 15856 6412 17408 6440
rect 15090 6344 15424 6372
rect 15090 6341 15102 6344
rect 15044 6335 15102 6341
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 11931 6276 11989 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 11977 6273 11989 6276
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 12066 6264 12072 6316
rect 12124 6304 12130 6316
rect 12161 6307 12219 6313
rect 12161 6304 12173 6307
rect 12124 6276 12173 6304
rect 12124 6264 12130 6276
rect 12161 6273 12173 6276
rect 12207 6273 12219 6307
rect 12161 6267 12219 6273
rect 8260 6208 8708 6236
rect 8260 6196 8266 6208
rect 9214 6196 9220 6248
rect 9272 6196 9278 6248
rect 9582 6196 9588 6248
rect 9640 6196 9646 6248
rect 9858 6196 9864 6248
rect 9916 6196 9922 6248
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6205 10011 6239
rect 13648 6236 13676 6335
rect 15488 6304 15516 6400
rect 15565 6307 15623 6313
rect 15565 6304 15577 6307
rect 15488 6276 15577 6304
rect 15565 6273 15577 6276
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 9953 6199 10011 6205
rect 13004 6208 13676 6236
rect 8113 6171 8171 6177
rect 8113 6137 8125 6171
rect 8159 6137 8171 6171
rect 8113 6131 8171 6137
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 9968 6168 9996 6199
rect 12158 6168 12164 6180
rect 8352 6140 9996 6168
rect 10888 6140 12164 6168
rect 8352 6128 8358 6140
rect 9582 6100 9588 6112
rect 7852 6072 9588 6100
rect 9582 6060 9588 6072
rect 9640 6100 9646 6112
rect 10888 6100 10916 6140
rect 12158 6128 12164 6140
rect 12216 6128 12222 6180
rect 13004 6177 13032 6208
rect 15286 6196 15292 6248
rect 15344 6196 15350 6248
rect 15856 6245 15884 6412
rect 17402 6400 17408 6412
rect 17460 6440 17466 6452
rect 17770 6440 17776 6452
rect 17460 6412 17776 6440
rect 17460 6400 17466 6412
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 18049 6443 18107 6449
rect 18049 6440 18061 6443
rect 17920 6412 18061 6440
rect 17920 6400 17926 6412
rect 18049 6409 18061 6412
rect 18095 6409 18107 6443
rect 18049 6403 18107 6409
rect 19521 6443 19579 6449
rect 19521 6409 19533 6443
rect 19567 6440 19579 6443
rect 19886 6440 19892 6452
rect 19567 6412 19892 6440
rect 19567 6409 19579 6412
rect 19521 6403 19579 6409
rect 19886 6400 19892 6412
rect 19944 6400 19950 6452
rect 19978 6372 19984 6384
rect 16684 6344 17908 6372
rect 16684 6313 16712 6344
rect 17880 6316 17908 6344
rect 18156 6344 19984 6372
rect 16669 6307 16727 6313
rect 16669 6273 16681 6307
rect 16715 6273 16727 6307
rect 16925 6307 16983 6313
rect 16925 6304 16937 6307
rect 16669 6267 16727 6273
rect 16776 6276 16937 6304
rect 15841 6239 15899 6245
rect 15841 6236 15853 6239
rect 15488 6208 15853 6236
rect 12989 6171 13047 6177
rect 12989 6137 13001 6171
rect 13035 6137 13047 6171
rect 12989 6131 13047 6137
rect 13262 6128 13268 6180
rect 13320 6128 13326 6180
rect 15488 6112 15516 6208
rect 15841 6205 15853 6208
rect 15887 6205 15899 6239
rect 15841 6199 15899 6205
rect 16022 6196 16028 6248
rect 16080 6236 16086 6248
rect 16776 6236 16804 6276
rect 16925 6273 16937 6276
rect 16971 6273 16983 6307
rect 16925 6267 16983 6273
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 18156 6313 18184 6344
rect 18141 6307 18199 6313
rect 18141 6304 18153 6307
rect 17920 6276 18153 6304
rect 17920 6264 17926 6276
rect 18141 6273 18153 6276
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 18408 6307 18466 6313
rect 18408 6273 18420 6307
rect 18454 6304 18466 6307
rect 18782 6304 18788 6316
rect 18454 6276 18788 6304
rect 18454 6273 18466 6276
rect 18408 6267 18466 6273
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 19628 6313 19656 6344
rect 19978 6332 19984 6344
rect 20036 6372 20042 6384
rect 20530 6372 20536 6384
rect 20036 6344 20536 6372
rect 20036 6332 20042 6344
rect 20530 6332 20536 6344
rect 20588 6332 20594 6384
rect 19613 6307 19671 6313
rect 19613 6273 19625 6307
rect 19659 6273 19671 6307
rect 19613 6267 19671 6273
rect 19880 6307 19938 6313
rect 19880 6273 19892 6307
rect 19926 6304 19938 6307
rect 20254 6304 20260 6316
rect 19926 6276 20260 6304
rect 19926 6273 19938 6276
rect 19880 6267 19938 6273
rect 20254 6264 20260 6276
rect 20312 6264 20318 6316
rect 16080 6208 16804 6236
rect 16080 6196 16086 6208
rect 9640 6072 10916 6100
rect 9640 6060 9646 6072
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 11333 6103 11391 6109
rect 11333 6100 11345 6103
rect 11204 6072 11345 6100
rect 11204 6060 11210 6072
rect 11333 6069 11345 6072
rect 11379 6069 11391 6103
rect 11333 6063 11391 6069
rect 13078 6060 13084 6112
rect 13136 6060 13142 6112
rect 15470 6060 15476 6112
rect 15528 6060 15534 6112
rect 16482 6060 16488 6112
rect 16540 6060 16546 6112
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 18046 6100 18052 6112
rect 16908 6072 18052 6100
rect 16908 6060 16914 6072
rect 18046 6060 18052 6072
rect 18104 6100 18110 6112
rect 19334 6100 19340 6112
rect 18104 6072 19340 6100
rect 18104 6060 18110 6072
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 20622 6060 20628 6112
rect 20680 6100 20686 6112
rect 20993 6103 21051 6109
rect 20993 6100 21005 6103
rect 20680 6072 21005 6100
rect 20680 6060 20686 6072
rect 20993 6069 21005 6072
rect 21039 6100 21051 6103
rect 21174 6100 21180 6112
rect 21039 6072 21180 6100
rect 21039 6069 21051 6072
rect 20993 6063 21051 6069
rect 21174 6060 21180 6072
rect 21232 6060 21238 6112
rect 1104 6010 22264 6032
rect 1104 5958 3595 6010
rect 3647 5958 3659 6010
rect 3711 5958 3723 6010
rect 3775 5958 3787 6010
rect 3839 5958 3851 6010
rect 3903 5958 8885 6010
rect 8937 5958 8949 6010
rect 9001 5958 9013 6010
rect 9065 5958 9077 6010
rect 9129 5958 9141 6010
rect 9193 5958 14175 6010
rect 14227 5958 14239 6010
rect 14291 5958 14303 6010
rect 14355 5958 14367 6010
rect 14419 5958 14431 6010
rect 14483 5958 19465 6010
rect 19517 5958 19529 6010
rect 19581 5958 19593 6010
rect 19645 5958 19657 6010
rect 19709 5958 19721 6010
rect 19773 5958 22264 6010
rect 1104 5936 22264 5958
rect 3234 5856 3240 5908
rect 3292 5896 3298 5908
rect 6457 5899 6515 5905
rect 3292 5868 5396 5896
rect 3292 5856 3298 5868
rect 3970 5652 3976 5704
rect 4028 5692 4034 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 4028 5664 4077 5692
rect 4028 5652 4034 5664
rect 4065 5661 4077 5664
rect 4111 5692 4123 5695
rect 4154 5692 4160 5704
rect 4111 5664 4160 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4332 5627 4390 5633
rect 4332 5593 4344 5627
rect 4378 5624 4390 5627
rect 4614 5624 4620 5636
rect 4378 5596 4620 5624
rect 4378 5593 4390 5596
rect 4332 5587 4390 5593
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 5368 5624 5396 5868
rect 6457 5865 6469 5899
rect 6503 5865 6515 5899
rect 6457 5859 6515 5865
rect 6917 5899 6975 5905
rect 6917 5865 6929 5899
rect 6963 5896 6975 5899
rect 7558 5896 7564 5908
rect 6963 5868 7564 5896
rect 6963 5865 6975 5868
rect 6917 5859 6975 5865
rect 5445 5831 5503 5837
rect 5445 5797 5457 5831
rect 5491 5797 5503 5831
rect 5445 5791 5503 5797
rect 5460 5692 5488 5791
rect 6270 5788 6276 5840
rect 6328 5788 6334 5840
rect 6472 5828 6500 5859
rect 7558 5856 7564 5868
rect 7616 5896 7622 5908
rect 7616 5868 8524 5896
rect 7616 5856 7622 5868
rect 7282 5828 7288 5840
rect 6472 5800 7288 5828
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 8496 5760 8524 5868
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 8628 5868 8677 5896
rect 8628 5856 8634 5868
rect 8665 5865 8677 5868
rect 8711 5865 8723 5899
rect 8665 5859 8723 5865
rect 9398 5856 9404 5908
rect 9456 5856 9462 5908
rect 9766 5856 9772 5908
rect 9824 5896 9830 5908
rect 9950 5896 9956 5908
rect 9824 5868 9956 5896
rect 9824 5856 9830 5868
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 13078 5856 13084 5908
rect 13136 5856 13142 5908
rect 15470 5856 15476 5908
rect 15528 5856 15534 5908
rect 16022 5856 16028 5908
rect 16080 5856 16086 5908
rect 16482 5856 16488 5908
rect 16540 5856 16546 5908
rect 20254 5856 20260 5908
rect 20312 5856 20318 5908
rect 9416 5828 9444 5856
rect 9416 5800 9674 5828
rect 9214 5760 9220 5772
rect 5592 5732 7328 5760
rect 8496 5732 9220 5760
rect 5592 5720 5598 5732
rect 6089 5695 6147 5701
rect 6089 5692 6101 5695
rect 5460 5664 6101 5692
rect 6089 5661 6101 5664
rect 6135 5661 6147 5695
rect 6914 5692 6920 5704
rect 6089 5655 6147 5661
rect 6380 5664 6920 5692
rect 6104 5624 6132 5655
rect 6380 5624 6408 5664
rect 6454 5633 6460 5636
rect 5368 5596 6040 5624
rect 6104 5596 6408 5624
rect 6441 5627 6460 5633
rect 5537 5559 5595 5565
rect 5537 5525 5549 5559
rect 5583 5556 5595 5559
rect 5626 5556 5632 5568
rect 5583 5528 5632 5556
rect 5583 5525 5595 5528
rect 5537 5519 5595 5525
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 6012 5556 6040 5596
rect 6441 5593 6453 5627
rect 6441 5587 6460 5593
rect 6454 5584 6460 5587
rect 6512 5584 6518 5636
rect 6656 5633 6684 5664
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 7300 5692 7328 5732
rect 9214 5720 9220 5732
rect 9272 5760 9278 5772
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 9272 5732 9413 5760
rect 9272 5720 9278 5732
rect 9401 5729 9413 5732
rect 9447 5729 9459 5763
rect 9646 5760 9674 5800
rect 9646 5732 10541 5760
rect 9401 5723 9459 5729
rect 8294 5692 8300 5704
rect 7300 5664 8300 5692
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5692 8631 5695
rect 8662 5692 8668 5704
rect 8619 5664 8668 5692
rect 8619 5661 8631 5664
rect 8573 5655 8631 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 6641 5627 6699 5633
rect 6641 5593 6653 5627
rect 6687 5593 6699 5627
rect 6641 5587 6699 5593
rect 8018 5584 8024 5636
rect 8076 5633 8082 5636
rect 8076 5627 8110 5633
rect 8098 5593 8110 5627
rect 8076 5587 8110 5593
rect 8076 5584 8082 5587
rect 8662 5556 8668 5568
rect 6012 5528 8668 5556
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 8772 5556 8800 5655
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9585 5695 9643 5701
rect 9585 5692 9597 5695
rect 8904 5664 9597 5692
rect 8904 5652 8910 5664
rect 9232 5636 9260 5664
rect 9585 5661 9597 5664
rect 9631 5692 9643 5695
rect 9631 5664 9812 5692
rect 9631 5661 9643 5664
rect 9585 5655 9643 5661
rect 9214 5584 9220 5636
rect 9272 5584 9278 5636
rect 9306 5584 9312 5636
rect 9364 5624 9370 5636
rect 9674 5624 9680 5636
rect 9364 5596 9680 5624
rect 9364 5584 9370 5596
rect 9674 5584 9680 5596
rect 9732 5584 9738 5636
rect 9398 5556 9404 5568
rect 8772 5528 9404 5556
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 9784 5556 9812 5664
rect 9858 5652 9864 5704
rect 9916 5652 9922 5704
rect 10410 5652 10416 5704
rect 10468 5652 10474 5704
rect 10513 5692 10541 5732
rect 10594 5720 10600 5772
rect 10652 5720 10658 5772
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5729 11299 5763
rect 11241 5723 11299 5729
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 10513 5664 10701 5692
rect 10689 5661 10701 5664
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 11146 5652 11152 5704
rect 11204 5652 11210 5704
rect 11256 5692 11284 5723
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11256 5664 11805 5692
rect 11256 5556 11284 5664
rect 11793 5661 11805 5664
rect 11839 5692 11851 5695
rect 12066 5692 12072 5704
rect 11839 5664 12072 5692
rect 11839 5661 11851 5664
rect 11793 5655 11851 5661
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5692 12955 5695
rect 13096 5692 13124 5856
rect 16500 5769 16528 5856
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5729 16543 5763
rect 16485 5723 16543 5729
rect 19613 5763 19671 5769
rect 19613 5729 19625 5763
rect 19659 5760 19671 5763
rect 19886 5760 19892 5772
rect 19659 5732 19892 5760
rect 19659 5729 19671 5732
rect 19613 5723 19671 5729
rect 19886 5720 19892 5732
rect 19944 5720 19950 5772
rect 21174 5720 21180 5772
rect 21232 5720 21238 5772
rect 12943 5664 13124 5692
rect 12943 5661 12955 5664
rect 12897 5655 12955 5661
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 13722 5692 13728 5704
rect 13320 5664 13728 5692
rect 13320 5652 13326 5664
rect 13722 5652 13728 5664
rect 13780 5692 13786 5704
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13780 5664 14105 5692
rect 13780 5652 13786 5664
rect 14093 5661 14105 5664
rect 14139 5692 14151 5695
rect 15286 5692 15292 5704
rect 14139 5664 15292 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5692 15899 5695
rect 16117 5695 16175 5701
rect 16117 5692 16129 5695
rect 15887 5664 16129 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 16117 5661 16129 5664
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 16301 5695 16359 5701
rect 16301 5661 16313 5695
rect 16347 5692 16359 5695
rect 16850 5692 16856 5704
rect 16347 5664 16856 5692
rect 16347 5661 16359 5664
rect 16301 5655 16359 5661
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 18138 5652 18144 5704
rect 18196 5692 18202 5704
rect 18601 5695 18659 5701
rect 18601 5692 18613 5695
rect 18196 5664 18613 5692
rect 18196 5652 18202 5664
rect 18601 5661 18613 5664
rect 18647 5661 18659 5695
rect 18601 5655 18659 5661
rect 20441 5695 20499 5701
rect 20441 5661 20453 5695
rect 20487 5692 20499 5695
rect 20530 5692 20536 5704
rect 20487 5664 20536 5692
rect 20487 5661 20499 5664
rect 20441 5655 20499 5661
rect 20530 5652 20536 5664
rect 20588 5652 20594 5704
rect 12158 5584 12164 5636
rect 12216 5624 12222 5636
rect 12216 5596 12434 5624
rect 12216 5584 12222 5596
rect 9784 5528 11284 5556
rect 12406 5556 12434 5596
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 14338 5627 14396 5633
rect 14338 5624 14350 5627
rect 13872 5596 14350 5624
rect 13872 5584 13878 5596
rect 14338 5593 14350 5596
rect 14384 5593 14396 5627
rect 14338 5587 14396 5593
rect 12713 5559 12771 5565
rect 12713 5556 12725 5559
rect 12406 5528 12725 5556
rect 12713 5525 12725 5528
rect 12759 5525 12771 5559
rect 12713 5519 12771 5525
rect 18046 5516 18052 5568
rect 18104 5516 18110 5568
rect 19886 5516 19892 5568
rect 19944 5556 19950 5568
rect 20165 5559 20223 5565
rect 20165 5556 20177 5559
rect 19944 5528 20177 5556
rect 19944 5516 19950 5528
rect 20165 5525 20177 5528
rect 20211 5525 20223 5559
rect 20165 5519 20223 5525
rect 20622 5516 20628 5568
rect 20680 5516 20686 5568
rect 1104 5466 22264 5488
rect 1104 5414 4255 5466
rect 4307 5414 4319 5466
rect 4371 5414 4383 5466
rect 4435 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 9545 5466
rect 9597 5414 9609 5466
rect 9661 5414 9673 5466
rect 9725 5414 9737 5466
rect 9789 5414 9801 5466
rect 9853 5414 14835 5466
rect 14887 5414 14899 5466
rect 14951 5414 14963 5466
rect 15015 5414 15027 5466
rect 15079 5414 15091 5466
rect 15143 5414 20125 5466
rect 20177 5414 20189 5466
rect 20241 5414 20253 5466
rect 20305 5414 20317 5466
rect 20369 5414 20381 5466
rect 20433 5414 22264 5466
rect 1104 5392 22264 5414
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4614 5352 4620 5364
rect 4571 5324 4620 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 7558 5312 7564 5364
rect 7616 5352 7622 5364
rect 9861 5355 9919 5361
rect 7616 5324 7880 5352
rect 7616 5312 7622 5324
rect 5169 5287 5227 5293
rect 5169 5284 5181 5287
rect 4724 5256 5181 5284
rect 4724 5225 4752 5256
rect 5169 5253 5181 5256
rect 5215 5253 5227 5287
rect 5169 5247 5227 5253
rect 5276 5256 5856 5284
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 4890 5176 4896 5228
rect 4948 5176 4954 5228
rect 5074 5176 5080 5228
rect 5132 5176 5138 5228
rect 5276 5225 5304 5256
rect 5828 5228 5856 5256
rect 6914 5244 6920 5296
rect 6972 5244 6978 5296
rect 7745 5287 7803 5293
rect 7745 5284 7757 5287
rect 7116 5256 7757 5284
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 5626 5176 5632 5228
rect 5684 5176 5690 5228
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 6086 5216 6092 5228
rect 5868 5188 6092 5216
rect 5868 5176 5874 5188
rect 6086 5176 6092 5188
rect 6144 5176 6150 5228
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5148 5043 5151
rect 5644 5148 5672 5176
rect 5031 5120 5672 5148
rect 6932 5148 6960 5244
rect 7116 5228 7144 5256
rect 7745 5253 7757 5256
rect 7791 5253 7803 5287
rect 7745 5247 7803 5253
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5216 7067 5219
rect 7098 5216 7104 5228
rect 7055 5188 7104 5216
rect 7055 5185 7067 5188
rect 7009 5179 7067 5185
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 7466 5216 7472 5228
rect 7423 5188 7472 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 7208 5148 7236 5179
rect 6932 5120 7236 5148
rect 7300 5148 7328 5179
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 7852 5225 7880 5324
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 10594 5352 10600 5364
rect 9907 5324 10600 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 14642 5312 14648 5364
rect 14700 5352 14706 5364
rect 15289 5355 15347 5361
rect 15289 5352 15301 5355
rect 14700 5324 15301 5352
rect 14700 5312 14706 5324
rect 15289 5321 15301 5324
rect 15335 5321 15347 5355
rect 15289 5315 15347 5321
rect 19334 5312 19340 5364
rect 19392 5312 19398 5364
rect 19705 5355 19763 5361
rect 19705 5321 19717 5355
rect 19751 5352 19763 5355
rect 19978 5352 19984 5364
rect 19751 5324 19984 5352
rect 19751 5321 19763 5324
rect 19705 5315 19763 5321
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20441 5355 20499 5361
rect 20441 5321 20453 5355
rect 20487 5352 20499 5355
rect 20530 5352 20536 5364
rect 20487 5324 20536 5352
rect 20487 5321 20499 5324
rect 20441 5315 20499 5321
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 20714 5312 20720 5364
rect 20772 5312 20778 5364
rect 20901 5355 20959 5361
rect 20901 5321 20913 5355
rect 20947 5352 20959 5355
rect 21818 5352 21824 5364
rect 20947 5324 21824 5352
rect 20947 5321 20959 5324
rect 20901 5315 20959 5321
rect 21818 5312 21824 5324
rect 21876 5312 21882 5364
rect 14734 5244 14740 5296
rect 14792 5284 14798 5296
rect 18233 5287 18291 5293
rect 18233 5284 18245 5287
rect 14792 5256 18245 5284
rect 14792 5244 14798 5256
rect 18233 5253 18245 5256
rect 18279 5253 18291 5287
rect 19352 5284 19380 5312
rect 19352 5256 20300 5284
rect 18233 5247 18291 5253
rect 7837 5219 7895 5225
rect 7837 5185 7849 5219
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5216 8447 5219
rect 9306 5216 9312 5228
rect 8435 5188 9312 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5216 9827 5219
rect 9858 5216 9864 5228
rect 9815 5188 9864 5216
rect 9815 5185 9827 5188
rect 9769 5179 9827 5185
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5216 10011 5219
rect 10042 5216 10048 5228
rect 9999 5188 10048 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 16022 5176 16028 5228
rect 16080 5176 16086 5228
rect 16390 5176 16396 5228
rect 16448 5216 16454 5228
rect 17126 5216 17132 5228
rect 16448 5188 17132 5216
rect 16448 5176 16454 5188
rect 17126 5176 17132 5188
rect 17184 5216 17190 5228
rect 17773 5219 17831 5225
rect 17773 5216 17785 5219
rect 17184 5188 17785 5216
rect 17184 5176 17190 5188
rect 17773 5185 17785 5188
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 17957 5219 18015 5225
rect 17957 5185 17969 5219
rect 18003 5216 18015 5219
rect 18046 5216 18052 5228
rect 18003 5188 18052 5216
rect 18003 5185 18015 5188
rect 17957 5179 18015 5185
rect 18046 5176 18052 5188
rect 18104 5176 18110 5228
rect 19886 5176 19892 5228
rect 19944 5216 19950 5228
rect 20272 5225 20300 5256
rect 20073 5219 20131 5225
rect 20073 5216 20085 5219
rect 19944 5188 20085 5216
rect 19944 5176 19950 5188
rect 20073 5185 20085 5188
rect 20119 5185 20131 5219
rect 20073 5179 20131 5185
rect 20257 5219 20315 5225
rect 20257 5185 20269 5219
rect 20303 5185 20315 5219
rect 20257 5179 20315 5185
rect 20622 5176 20628 5228
rect 20680 5176 20686 5228
rect 20732 5225 20760 5312
rect 20717 5219 20775 5225
rect 20717 5185 20729 5219
rect 20763 5185 20775 5219
rect 20717 5179 20775 5185
rect 7742 5148 7748 5160
rect 7300 5120 7748 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 7742 5108 7748 5120
rect 7800 5148 7806 5160
rect 8297 5151 8355 5157
rect 8297 5148 8309 5151
rect 7800 5120 8309 5148
rect 7800 5108 7806 5120
rect 8297 5117 8309 5120
rect 8343 5117 8355 5151
rect 8297 5111 8355 5117
rect 16298 5108 16304 5160
rect 16356 5108 16362 5160
rect 2746 5052 7696 5080
rect 1854 4972 1860 5024
rect 1912 5012 1918 5024
rect 2746 5012 2774 5052
rect 7668 5024 7696 5052
rect 1912 4984 2774 5012
rect 1912 4972 1918 4984
rect 7558 4972 7564 5024
rect 7616 4972 7622 5024
rect 7650 4972 7656 5024
rect 7708 4972 7714 5024
rect 12894 4972 12900 5024
rect 12952 5012 12958 5024
rect 13262 5012 13268 5024
rect 12952 4984 13268 5012
rect 12952 4972 12958 4984
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 16408 5012 16436 5176
rect 15436 4984 16436 5012
rect 15436 4972 15442 4984
rect 17218 4972 17224 5024
rect 17276 5012 17282 5024
rect 17589 5015 17647 5021
rect 17589 5012 17601 5015
rect 17276 4984 17601 5012
rect 17276 4972 17282 4984
rect 17589 4981 17601 4984
rect 17635 4981 17647 5015
rect 17589 4975 17647 4981
rect 1104 4922 22264 4944
rect 1104 4870 3595 4922
rect 3647 4870 3659 4922
rect 3711 4870 3723 4922
rect 3775 4870 3787 4922
rect 3839 4870 3851 4922
rect 3903 4870 8885 4922
rect 8937 4870 8949 4922
rect 9001 4870 9013 4922
rect 9065 4870 9077 4922
rect 9129 4870 9141 4922
rect 9193 4870 14175 4922
rect 14227 4870 14239 4922
rect 14291 4870 14303 4922
rect 14355 4870 14367 4922
rect 14419 4870 14431 4922
rect 14483 4870 19465 4922
rect 19517 4870 19529 4922
rect 19581 4870 19593 4922
rect 19645 4870 19657 4922
rect 19709 4870 19721 4922
rect 19773 4870 22264 4922
rect 1104 4848 22264 4870
rect 6270 4808 6276 4820
rect 5552 4780 6276 4808
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 5074 4604 5080 4616
rect 4856 4576 5080 4604
rect 4856 4564 4862 4576
rect 5074 4564 5080 4576
rect 5132 4604 5138 4616
rect 5552 4613 5580 4780
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 7558 4768 7564 4820
rect 7616 4768 7622 4820
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 13722 4808 13728 4820
rect 7708 4780 13728 4808
rect 7708 4768 7714 4780
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 13814 4768 13820 4820
rect 13872 4768 13878 4820
rect 15746 4768 15752 4820
rect 15804 4768 15810 4820
rect 16022 4768 16028 4820
rect 16080 4768 16086 4820
rect 16117 4811 16175 4817
rect 16117 4777 16129 4811
rect 16163 4808 16175 4811
rect 16298 4808 16304 4820
rect 16163 4780 16304 4808
rect 16163 4777 16175 4780
rect 16117 4771 16175 4777
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 17218 4808 17224 4820
rect 16776 4780 17224 4808
rect 7466 4700 7472 4752
rect 7524 4700 7530 4752
rect 5902 4672 5908 4684
rect 5736 4644 5908 4672
rect 5736 4613 5764 4644
rect 5902 4632 5908 4644
rect 5960 4672 5966 4684
rect 7484 4672 7512 4700
rect 7576 4681 7604 4768
rect 7742 4700 7748 4752
rect 7800 4700 7806 4752
rect 11698 4700 11704 4752
rect 11756 4740 11762 4752
rect 15764 4740 15792 4768
rect 11756 4712 15792 4740
rect 16040 4740 16068 4768
rect 16209 4743 16267 4749
rect 16209 4740 16221 4743
rect 16040 4712 16221 4740
rect 11756 4700 11762 4712
rect 5960 4644 7512 4672
rect 7561 4675 7619 4681
rect 5960 4632 5966 4644
rect 7561 4641 7573 4675
rect 7607 4641 7619 4675
rect 7561 4635 7619 4641
rect 7650 4632 7656 4684
rect 7708 4632 7714 4684
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 5132 4576 5549 4604
rect 5132 4564 5138 4576
rect 5537 4573 5549 4576
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 5350 4496 5356 4548
rect 5408 4536 5414 4548
rect 6012 4536 6040 4567
rect 6086 4564 6092 4616
rect 6144 4604 6150 4616
rect 6181 4607 6239 4613
rect 6181 4604 6193 4607
rect 6144 4576 6193 4604
rect 6144 4564 6150 4576
rect 6181 4573 6193 4576
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 7282 4564 7288 4616
rect 7340 4564 7346 4616
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 7432 4576 7481 4604
rect 7432 4564 7438 4576
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 7760 4604 7788 4700
rect 13280 4613 13308 4712
rect 14829 4675 14887 4681
rect 14829 4641 14841 4675
rect 14875 4672 14887 4675
rect 15194 4672 15200 4684
rect 14875 4644 15200 4672
rect 14875 4641 14887 4644
rect 14829 4635 14887 4641
rect 15194 4632 15200 4644
rect 15252 4632 15258 4684
rect 7837 4607 7895 4613
rect 7837 4604 7849 4607
rect 7760 4576 7849 4604
rect 7469 4567 7527 4573
rect 7837 4573 7849 4576
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 13265 4607 13323 4613
rect 13265 4573 13277 4607
rect 13311 4573 13323 4607
rect 13265 4567 13323 4573
rect 13630 4564 13636 4616
rect 13688 4564 13694 4616
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4604 15071 4607
rect 15378 4604 15384 4616
rect 15059 4576 15384 4604
rect 15059 4573 15071 4576
rect 15013 4567 15071 4573
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 15473 4607 15531 4613
rect 15473 4573 15485 4607
rect 15519 4573 15531 4607
rect 15473 4567 15531 4573
rect 5408 4508 6040 4536
rect 15488 4536 15516 4567
rect 15654 4564 15660 4616
rect 15712 4564 15718 4616
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16040 4604 16068 4712
rect 16209 4709 16221 4712
rect 16255 4709 16267 4743
rect 16209 4703 16267 4709
rect 15979 4576 16068 4604
rect 16393 4607 16451 4613
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 16393 4573 16405 4607
rect 16439 4604 16451 4607
rect 16666 4604 16672 4616
rect 16439 4576 16672 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 16776 4613 16804 4780
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 16761 4607 16819 4613
rect 16761 4573 16773 4607
rect 16807 4573 16819 4607
rect 16761 4567 16819 4573
rect 17037 4607 17095 4613
rect 17037 4573 17049 4607
rect 17083 4604 17095 4607
rect 17862 4604 17868 4616
rect 17083 4576 17868 4604
rect 17083 4573 17095 4576
rect 17037 4567 17095 4573
rect 17862 4564 17868 4576
rect 17920 4564 17926 4616
rect 18506 4564 18512 4616
rect 18564 4564 18570 4616
rect 16850 4536 16856 4548
rect 15488 4508 16856 4536
rect 5408 4496 5414 4508
rect 16850 4496 16856 4508
rect 16908 4496 16914 4548
rect 17282 4539 17340 4545
rect 17282 4536 17294 4539
rect 16960 4508 17294 4536
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 6089 4471 6147 4477
rect 6089 4468 6101 4471
rect 5684 4440 6101 4468
rect 5684 4428 5690 4440
rect 6089 4437 6101 4440
rect 6135 4437 6147 4471
rect 6089 4431 6147 4437
rect 8021 4471 8079 4477
rect 8021 4437 8033 4471
rect 8067 4468 8079 4471
rect 8110 4468 8116 4480
rect 8067 4440 8116 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 13449 4471 13507 4477
rect 13449 4437 13461 4471
rect 13495 4468 13507 4471
rect 13722 4468 13728 4480
rect 13495 4440 13728 4468
rect 13495 4437 13507 4440
rect 13449 4431 13507 4437
rect 13722 4428 13728 4440
rect 13780 4428 13786 4480
rect 15197 4471 15255 4477
rect 15197 4437 15209 4471
rect 15243 4468 15255 4471
rect 16206 4468 16212 4480
rect 15243 4440 16212 4468
rect 15243 4437 15255 4440
rect 15197 4431 15255 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 16960 4477 16988 4508
rect 17282 4505 17294 4508
rect 17328 4505 17340 4539
rect 17282 4499 17340 4505
rect 16945 4471 17003 4477
rect 16945 4437 16957 4471
rect 16991 4437 17003 4471
rect 16945 4431 17003 4437
rect 18414 4428 18420 4480
rect 18472 4428 18478 4480
rect 18690 4428 18696 4480
rect 18748 4428 18754 4480
rect 1104 4378 22264 4400
rect 1104 4326 4255 4378
rect 4307 4326 4319 4378
rect 4371 4326 4383 4378
rect 4435 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 9545 4378
rect 9597 4326 9609 4378
rect 9661 4326 9673 4378
rect 9725 4326 9737 4378
rect 9789 4326 9801 4378
rect 9853 4326 14835 4378
rect 14887 4326 14899 4378
rect 14951 4326 14963 4378
rect 15015 4326 15027 4378
rect 15079 4326 15091 4378
rect 15143 4326 20125 4378
rect 20177 4326 20189 4378
rect 20241 4326 20253 4378
rect 20305 4326 20317 4378
rect 20369 4326 20381 4378
rect 20433 4326 22264 4378
rect 1104 4304 22264 4326
rect 11698 4264 11704 4276
rect 10980 4236 11704 4264
rect 7926 4156 7932 4208
rect 7984 4196 7990 4208
rect 9766 4196 9772 4208
rect 7984 4168 8616 4196
rect 7984 4156 7990 4168
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 4663 4100 5120 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 4798 4020 4804 4072
rect 4856 4020 4862 4072
rect 4893 4063 4951 4069
rect 4893 4029 4905 4063
rect 4939 4029 4951 4063
rect 5092 4060 5120 4100
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 5350 4088 5356 4140
rect 5408 4088 5414 4140
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 5491 4100 6377 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 6365 4091 6423 4097
rect 6840 4100 7389 4128
rect 5626 4060 5632 4072
rect 5092 4032 5632 4060
rect 4893 4023 4951 4029
rect 4908 3992 4936 4023
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 5902 4020 5908 4072
rect 5960 4060 5966 4072
rect 6089 4063 6147 4069
rect 6089 4060 6101 4063
rect 5960 4032 6101 4060
rect 5960 4020 5966 4032
rect 6089 4029 6101 4032
rect 6135 4029 6147 4063
rect 6089 4023 6147 4029
rect 5537 3995 5595 4001
rect 5537 3992 5549 3995
rect 4908 3964 5549 3992
rect 5537 3961 5549 3964
rect 5583 3961 5595 3995
rect 5537 3955 5595 3961
rect 6840 3936 6868 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 8018 4088 8024 4140
rect 8076 4128 8082 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 8076 4100 8125 4128
rect 8076 4088 8082 4100
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 6917 4063 6975 4069
rect 6917 4029 6929 4063
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 6932 3936 6960 4023
rect 8021 3995 8079 4001
rect 8021 3961 8033 3995
rect 8067 3992 8079 3995
rect 8220 3992 8248 4091
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 8067 3964 8524 3992
rect 8067 3961 8079 3964
rect 8021 3955 8079 3961
rect 8496 3936 8524 3964
rect 4433 3927 4491 3933
rect 4433 3893 4445 3927
rect 4479 3924 4491 3927
rect 4614 3924 4620 3936
rect 4479 3896 4620 3924
rect 4479 3893 4491 3896
rect 4433 3887 4491 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3924 5043 3927
rect 5074 3924 5080 3936
rect 5031 3896 5080 3924
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 6822 3884 6828 3936
rect 6880 3884 6886 3936
rect 6914 3884 6920 3936
rect 6972 3884 6978 3936
rect 8202 3884 8208 3936
rect 8260 3924 8266 3936
rect 8389 3927 8447 3933
rect 8389 3924 8401 3927
rect 8260 3896 8401 3924
rect 8260 3884 8266 3896
rect 8389 3893 8401 3896
rect 8435 3893 8447 3927
rect 8389 3887 8447 3893
rect 8478 3884 8484 3936
rect 8536 3884 8542 3936
rect 8588 3924 8616 4168
rect 9140 4168 9772 4196
rect 8662 4088 8668 4140
rect 8720 4128 8726 4140
rect 9140 4128 9168 4168
rect 9766 4156 9772 4168
rect 9824 4156 9830 4208
rect 10980 4205 11008 4236
rect 11698 4224 11704 4236
rect 11756 4224 11762 4276
rect 15194 4224 15200 4276
rect 15252 4224 15258 4276
rect 15378 4224 15384 4276
rect 15436 4224 15442 4276
rect 16666 4224 16672 4276
rect 16724 4224 16730 4276
rect 17589 4267 17647 4273
rect 17589 4233 17601 4267
rect 17635 4264 17647 4267
rect 17678 4264 17684 4276
rect 17635 4236 17684 4264
rect 17635 4233 17647 4236
rect 17589 4227 17647 4233
rect 17678 4224 17684 4236
rect 17736 4224 17742 4276
rect 17773 4267 17831 4273
rect 17773 4233 17785 4267
rect 17819 4264 17831 4267
rect 17862 4264 17868 4276
rect 17819 4236 17868 4264
rect 17819 4233 17831 4236
rect 17773 4227 17831 4233
rect 17862 4224 17868 4236
rect 17920 4264 17926 4276
rect 18414 4264 18420 4276
rect 17920 4236 18420 4264
rect 17920 4224 17926 4236
rect 18414 4224 18420 4236
rect 18472 4224 18478 4276
rect 19978 4224 19984 4276
rect 20036 4224 20042 4276
rect 10965 4199 11023 4205
rect 10965 4165 10977 4199
rect 11011 4165 11023 4199
rect 10965 4159 11023 4165
rect 11181 4199 11239 4205
rect 11181 4165 11193 4199
rect 11227 4196 11239 4199
rect 12618 4196 12624 4208
rect 11227 4168 12624 4196
rect 11227 4165 11239 4168
rect 11181 4159 11239 4165
rect 12618 4156 12624 4168
rect 12676 4156 12682 4208
rect 13722 4156 13728 4208
rect 13780 4196 13786 4208
rect 15396 4196 15424 4224
rect 13780 4168 15424 4196
rect 15933 4199 15991 4205
rect 13780 4156 13786 4168
rect 8720 4100 9168 4128
rect 8720 4088 8726 4100
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 9272 4100 9413 4128
rect 9272 4088 9278 4100
rect 9401 4097 9413 4100
rect 9447 4097 9459 4131
rect 9401 4091 9459 4097
rect 9582 4088 9588 4140
rect 9640 4088 9646 4140
rect 9953 4131 10011 4137
rect 9953 4128 9965 4131
rect 9692 4100 9965 4128
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4060 9551 4063
rect 9692 4060 9720 4100
rect 9953 4097 9965 4100
rect 9999 4097 10011 4131
rect 11517 4131 11575 4137
rect 11517 4126 11529 4131
rect 9953 4091 10011 4097
rect 11440 4098 11529 4126
rect 9539 4032 9720 4060
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 9600 4004 9628 4032
rect 9766 4020 9772 4072
rect 9824 4020 9830 4072
rect 11440 4060 11468 4098
rect 11517 4097 11529 4098
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 14016 4137 14044 4168
rect 15933 4165 15945 4199
rect 15979 4165 15991 4199
rect 15933 4159 15991 4165
rect 12906 4131 12964 4137
rect 12906 4128 12918 4131
rect 11756 4100 12918 4128
rect 11756 4088 11762 4100
rect 12906 4097 12918 4100
rect 12952 4097 12964 4131
rect 12906 4091 12964 4097
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13311 4100 13829 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4128 15899 4131
rect 15948 4128 15976 4159
rect 16114 4156 16120 4208
rect 16172 4205 16178 4208
rect 16172 4199 16191 4205
rect 16179 4165 16191 4199
rect 16172 4159 16191 4165
rect 16172 4156 16178 4159
rect 16482 4156 16488 4208
rect 16540 4156 16546 4208
rect 16821 4199 16879 4205
rect 16821 4196 16833 4199
rect 16592 4168 16833 4196
rect 16500 4128 16528 4156
rect 15887 4100 16528 4128
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 11348 4032 11468 4060
rect 13173 4063 13231 4069
rect 9582 3952 9588 4004
rect 9640 3952 9646 4004
rect 11348 4001 11376 4032
rect 13173 4029 13185 4063
rect 13219 4029 13231 4063
rect 13173 4023 13231 4029
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4060 14243 4063
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 14231 4032 14289 4060
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 14277 4023 14335 4029
rect 14752 4032 14841 4060
rect 11333 3995 11391 4001
rect 9968 3964 11284 3992
rect 9968 3924 9996 3964
rect 8588 3896 9996 3924
rect 10137 3927 10195 3933
rect 10137 3893 10149 3927
rect 10183 3924 10195 3927
rect 10686 3924 10692 3936
rect 10183 3896 10692 3924
rect 10183 3893 10195 3896
rect 10137 3887 10195 3893
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 11149 3927 11207 3933
rect 11149 3924 11161 3927
rect 11112 3896 11161 3924
rect 11112 3884 11118 3896
rect 11149 3893 11161 3896
rect 11195 3893 11207 3927
rect 11256 3924 11284 3964
rect 11333 3961 11345 3995
rect 11379 3961 11391 3995
rect 11333 3955 11391 3961
rect 11698 3952 11704 4004
rect 11756 3952 11762 4004
rect 11790 3924 11796 3936
rect 11256 3896 11796 3924
rect 11149 3887 11207 3893
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 13188 3924 13216 4023
rect 14752 3936 14780 4032
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 16301 3995 16359 4001
rect 16301 3961 16313 3995
rect 16347 3992 16359 3995
rect 16592 3992 16620 4168
rect 16821 4165 16833 4168
rect 16867 4165 16879 4199
rect 16821 4159 16879 4165
rect 17034 4156 17040 4208
rect 17092 4156 17098 4208
rect 18690 4156 18696 4208
rect 18748 4196 18754 4208
rect 19162 4199 19220 4205
rect 19162 4196 19174 4199
rect 18748 4168 19174 4196
rect 18748 4156 18754 4168
rect 19162 4165 19174 4168
rect 19208 4165 19220 4199
rect 19162 4159 19220 4165
rect 19996 4196 20024 4224
rect 19996 4168 20760 4196
rect 17681 4131 17739 4137
rect 17681 4097 17693 4131
rect 17727 4097 17739 4131
rect 17681 4091 17739 4097
rect 16347 3964 16620 3992
rect 16347 3961 16359 3964
rect 16301 3955 16359 3961
rect 12952 3896 13216 3924
rect 12952 3884 12958 3896
rect 13446 3884 13452 3936
rect 13504 3884 13510 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 16117 3927 16175 3933
rect 16117 3924 16129 3927
rect 14792 3896 16129 3924
rect 14792 3884 14798 3896
rect 16117 3893 16129 3896
rect 16163 3924 16175 3927
rect 16574 3924 16580 3936
rect 16163 3896 16580 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 16853 3927 16911 3933
rect 16853 3893 16865 3927
rect 16899 3924 16911 3927
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 16899 3896 17417 3924
rect 16899 3893 16911 3896
rect 16853 3887 16911 3893
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 17696 3924 17724 4091
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 19392 4100 19441 4128
rect 19392 4088 19398 4100
rect 19429 4097 19441 4100
rect 19475 4128 19487 4131
rect 19996 4128 20024 4168
rect 19475 4100 20024 4128
rect 19475 4097 19487 4100
rect 19429 4091 19487 4097
rect 20162 4088 20168 4140
rect 20220 4128 20226 4140
rect 20634 4131 20692 4137
rect 20634 4128 20646 4131
rect 20220 4100 20646 4128
rect 20220 4088 20226 4100
rect 20634 4097 20646 4100
rect 20680 4097 20692 4131
rect 20732 4128 20760 4168
rect 20901 4131 20959 4137
rect 20901 4128 20913 4131
rect 20732 4100 20913 4128
rect 20634 4091 20692 4097
rect 20901 4097 20913 4100
rect 20947 4097 20959 4131
rect 20901 4091 20959 4097
rect 17957 4063 18015 4069
rect 17957 4029 17969 4063
rect 18003 4060 18015 4063
rect 18046 4060 18052 4072
rect 18003 4032 18052 4060
rect 18003 4029 18015 4032
rect 17957 4023 18015 4029
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 17770 3924 17776 3936
rect 17696 3896 17776 3924
rect 17405 3887 17463 3893
rect 17770 3884 17776 3896
rect 17828 3924 17834 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 17828 3896 18061 3924
rect 17828 3884 17834 3896
rect 18049 3893 18061 3896
rect 18095 3924 18107 3927
rect 18138 3924 18144 3936
rect 18095 3896 18144 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 19521 3927 19579 3933
rect 19521 3893 19533 3927
rect 19567 3924 19579 3927
rect 19794 3924 19800 3936
rect 19567 3896 19800 3924
rect 19567 3893 19579 3896
rect 19521 3887 19579 3893
rect 19794 3884 19800 3896
rect 19852 3884 19858 3936
rect 1104 3834 22264 3856
rect 1104 3782 3595 3834
rect 3647 3782 3659 3834
rect 3711 3782 3723 3834
rect 3775 3782 3787 3834
rect 3839 3782 3851 3834
rect 3903 3782 8885 3834
rect 8937 3782 8949 3834
rect 9001 3782 9013 3834
rect 9065 3782 9077 3834
rect 9129 3782 9141 3834
rect 9193 3782 14175 3834
rect 14227 3782 14239 3834
rect 14291 3782 14303 3834
rect 14355 3782 14367 3834
rect 14419 3782 14431 3834
rect 14483 3782 19465 3834
rect 19517 3782 19529 3834
rect 19581 3782 19593 3834
rect 19645 3782 19657 3834
rect 19709 3782 19721 3834
rect 19773 3782 22264 3834
rect 1104 3760 22264 3782
rect 7193 3723 7251 3729
rect 7193 3689 7205 3723
rect 7239 3720 7251 3723
rect 7282 3720 7288 3732
rect 7239 3692 7288 3720
rect 7239 3689 7251 3692
rect 7193 3683 7251 3689
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 7377 3723 7435 3729
rect 7377 3689 7389 3723
rect 7423 3689 7435 3723
rect 7377 3683 7435 3689
rect 6365 3655 6423 3661
rect 6365 3621 6377 3655
rect 6411 3652 6423 3655
rect 6914 3652 6920 3664
rect 6411 3624 6920 3652
rect 6411 3621 6423 3624
rect 6365 3615 6423 3621
rect 6914 3612 6920 3624
rect 6972 3652 6978 3664
rect 7009 3655 7067 3661
rect 7009 3652 7021 3655
rect 6972 3624 7021 3652
rect 6972 3612 6978 3624
rect 7009 3621 7021 3624
rect 7055 3652 7067 3655
rect 7392 3652 7420 3683
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 8665 3723 8723 3729
rect 8665 3720 8677 3723
rect 8444 3692 8677 3720
rect 8444 3680 8450 3692
rect 8665 3689 8677 3692
rect 8711 3689 8723 3723
rect 8665 3683 8723 3689
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9766 3720 9772 3732
rect 9539 3692 9772 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 7055 3624 7420 3652
rect 7055 3621 7067 3624
rect 7009 3615 7067 3621
rect 8018 3612 8024 3664
rect 8076 3652 8082 3664
rect 8573 3655 8631 3661
rect 8573 3652 8585 3655
rect 8076 3624 8585 3652
rect 8076 3612 8082 3624
rect 8573 3621 8585 3624
rect 8619 3621 8631 3655
rect 8573 3615 8631 3621
rect 9582 3612 9588 3664
rect 9640 3612 9646 3664
rect 7101 3587 7159 3593
rect 7101 3553 7113 3587
rect 7147 3584 7159 3587
rect 8297 3587 8355 3593
rect 7147 3556 8064 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3516 5043 3519
rect 5534 3516 5540 3528
rect 5031 3488 5540 3516
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3516 6699 3519
rect 7653 3519 7711 3525
rect 7653 3516 7665 3519
rect 6687 3488 7665 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 7653 3485 7665 3488
rect 7699 3516 7711 3519
rect 7926 3516 7932 3528
rect 7699 3488 7932 3516
rect 7699 3485 7711 3488
rect 7653 3479 7711 3485
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8036 3525 8064 3556
rect 8297 3553 8309 3587
rect 8343 3553 8355 3587
rect 8297 3547 8355 3553
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 8110 3476 8116 3528
rect 8168 3476 8174 3528
rect 5074 3408 5080 3460
rect 5132 3448 5138 3460
rect 5230 3451 5288 3457
rect 5230 3448 5242 3451
rect 5132 3420 5242 3448
rect 5132 3408 5138 3420
rect 5230 3417 5242 3420
rect 5276 3417 5288 3451
rect 5230 3411 5288 3417
rect 6822 3408 6828 3460
rect 6880 3448 6886 3460
rect 8312 3448 8340 3547
rect 8662 3544 8668 3596
rect 8720 3584 8726 3596
rect 8757 3587 8815 3593
rect 8757 3584 8769 3587
rect 8720 3556 8769 3584
rect 8720 3544 8726 3556
rect 8757 3553 8769 3556
rect 8803 3553 8815 3587
rect 8757 3547 8815 3553
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 6880 3420 8340 3448
rect 8404 3448 8432 3479
rect 8478 3476 8484 3528
rect 8536 3476 8542 3528
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3516 9183 3519
rect 9214 3516 9220 3528
rect 9171 3488 9220 3516
rect 9171 3485 9183 3488
rect 9125 3479 9183 3485
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9600 3525 9628 3612
rect 9692 3525 9720 3692
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 9953 3723 10011 3729
rect 9953 3689 9965 3723
rect 9999 3689 10011 3723
rect 11238 3720 11244 3732
rect 9953 3683 10011 3689
rect 10520 3692 11244 3720
rect 9968 3652 9996 3683
rect 10520 3661 10548 3692
rect 11238 3680 11244 3692
rect 11296 3720 11302 3732
rect 11296 3692 12388 3720
rect 11296 3680 11302 3692
rect 10321 3655 10379 3661
rect 10321 3652 10333 3655
rect 9968 3624 10333 3652
rect 10321 3621 10333 3624
rect 10367 3621 10379 3655
rect 10321 3615 10379 3621
rect 10505 3655 10563 3661
rect 10505 3621 10517 3655
rect 10551 3621 10563 3655
rect 10505 3615 10563 3621
rect 10686 3612 10692 3664
rect 10744 3612 10750 3664
rect 12360 3652 12388 3692
rect 12434 3680 12440 3732
rect 12492 3680 12498 3732
rect 12618 3680 12624 3732
rect 12676 3720 12682 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 12676 3692 12909 3720
rect 12676 3680 12682 3692
rect 12897 3689 12909 3692
rect 12943 3689 12955 3723
rect 12897 3683 12955 3689
rect 13357 3723 13415 3729
rect 13357 3689 13369 3723
rect 13403 3720 13415 3723
rect 13630 3720 13636 3732
rect 13403 3692 13636 3720
rect 13403 3689 13415 3692
rect 13357 3683 13415 3689
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 15654 3680 15660 3732
rect 15712 3720 15718 3732
rect 16301 3723 16359 3729
rect 16301 3720 16313 3723
rect 15712 3692 16313 3720
rect 15712 3680 15718 3692
rect 16301 3689 16313 3692
rect 16347 3689 16359 3723
rect 16301 3683 16359 3689
rect 16482 3680 16488 3732
rect 16540 3680 16546 3732
rect 16850 3680 16856 3732
rect 16908 3720 16914 3732
rect 17405 3723 17463 3729
rect 17405 3720 17417 3723
rect 16908 3692 17417 3720
rect 16908 3680 16914 3692
rect 17405 3689 17417 3692
rect 17451 3689 17463 3723
rect 17405 3683 17463 3689
rect 17862 3680 17868 3732
rect 17920 3720 17926 3732
rect 17920 3692 18092 3720
rect 17920 3680 17926 3692
rect 15473 3655 15531 3661
rect 12360 3624 12664 3652
rect 12529 3587 12587 3593
rect 12529 3584 12541 3587
rect 10796 3556 12112 3584
rect 9585 3519 9643 3525
rect 9585 3485 9597 3519
rect 9631 3485 9643 3519
rect 9585 3479 9643 3485
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3485 9735 3519
rect 9677 3479 9735 3485
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3516 10103 3519
rect 10502 3516 10508 3528
rect 10091 3488 10508 3516
rect 10091 3485 10103 3488
rect 10045 3479 10103 3485
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 10594 3476 10600 3528
rect 10652 3476 10658 3528
rect 10796 3525 10824 3556
rect 12084 3528 12112 3556
rect 12268 3556 12541 3584
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3485 10839 3519
rect 10781 3479 10839 3485
rect 10870 3476 10876 3528
rect 10928 3516 10934 3528
rect 11057 3519 11115 3525
rect 11057 3516 11069 3519
rect 10928 3488 11069 3516
rect 10928 3476 10934 3488
rect 11057 3485 11069 3488
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 11204 3488 11621 3516
rect 11204 3476 11210 3488
rect 11609 3485 11621 3488
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 11977 3519 12035 3525
rect 11977 3485 11989 3519
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 9309 3451 9367 3457
rect 8404 3420 8616 3448
rect 6880 3408 6886 3420
rect 7837 3383 7895 3389
rect 7837 3349 7849 3383
rect 7883 3380 7895 3383
rect 8478 3380 8484 3392
rect 7883 3352 8484 3380
rect 7883 3349 7895 3352
rect 7837 3343 7895 3349
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 8588 3380 8616 3420
rect 9309 3417 9321 3451
rect 9355 3417 9367 3451
rect 11793 3451 11851 3457
rect 11793 3448 11805 3451
rect 9309 3411 9367 3417
rect 9784 3420 11805 3448
rect 9324 3380 9352 3411
rect 9398 3380 9404 3392
rect 8588 3352 9404 3380
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 9784 3389 9812 3420
rect 11793 3417 11805 3420
rect 11839 3417 11851 3451
rect 11793 3411 11851 3417
rect 11992 3448 12020 3479
rect 12066 3476 12072 3528
rect 12124 3476 12130 3528
rect 12158 3476 12164 3528
rect 12216 3516 12222 3528
rect 12268 3525 12296 3556
rect 12529 3553 12541 3556
rect 12575 3553 12587 3587
rect 12529 3547 12587 3553
rect 12253 3519 12311 3525
rect 12253 3516 12265 3519
rect 12216 3488 12265 3516
rect 12216 3476 12222 3488
rect 12253 3485 12265 3488
rect 12299 3485 12311 3519
rect 12253 3479 12311 3485
rect 12345 3519 12403 3525
rect 12345 3485 12357 3519
rect 12391 3516 12403 3519
rect 12636 3516 12664 3624
rect 15473 3621 15485 3655
rect 15519 3652 15531 3655
rect 16500 3652 16528 3680
rect 15519 3624 16528 3652
rect 17313 3655 17371 3661
rect 15519 3621 15531 3624
rect 15473 3615 15531 3621
rect 17313 3621 17325 3655
rect 17359 3652 17371 3655
rect 17954 3652 17960 3664
rect 17359 3624 17960 3652
rect 17359 3621 17371 3624
rect 17313 3615 17371 3621
rect 17954 3612 17960 3624
rect 18012 3612 18018 3664
rect 12894 3544 12900 3596
rect 12952 3584 12958 3596
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 12952 3556 14105 3584
rect 12952 3544 12958 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 16114 3544 16120 3596
rect 16172 3584 16178 3596
rect 16390 3584 16396 3596
rect 16172 3556 16396 3584
rect 16172 3544 16178 3556
rect 16390 3544 16396 3556
rect 16448 3584 16454 3596
rect 16945 3587 17003 3593
rect 16448 3556 16804 3584
rect 16448 3544 16454 3556
rect 12713 3519 12771 3525
rect 12713 3516 12725 3519
rect 12391 3488 12725 3516
rect 12391 3485 12403 3488
rect 12345 3479 12403 3485
rect 12713 3485 12725 3488
rect 12759 3485 12771 3519
rect 12713 3479 12771 3485
rect 12986 3476 12992 3528
rect 13044 3476 13050 3528
rect 13170 3476 13176 3528
rect 13228 3476 13234 3528
rect 13446 3476 13452 3528
rect 13504 3476 13510 3528
rect 13633 3519 13691 3525
rect 13633 3485 13645 3519
rect 13679 3516 13691 3519
rect 13722 3516 13728 3528
rect 13679 3488 13728 3516
rect 13679 3485 13691 3488
rect 13633 3479 13691 3485
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 13817 3519 13875 3525
rect 13817 3485 13829 3519
rect 13863 3516 13875 3519
rect 15565 3519 15623 3525
rect 15565 3516 15577 3519
rect 13863 3488 15577 3516
rect 13863 3485 13875 3488
rect 13817 3479 13875 3485
rect 15565 3485 15577 3488
rect 15611 3485 15623 3519
rect 15565 3479 15623 3485
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3485 16543 3519
rect 16485 3479 16543 3485
rect 12437 3451 12495 3457
rect 12437 3448 12449 3451
rect 11992 3420 12449 3448
rect 9769 3383 9827 3389
rect 9769 3349 9781 3383
rect 9815 3349 9827 3383
rect 9769 3343 9827 3349
rect 10042 3340 10048 3392
rect 10100 3340 10106 3392
rect 10410 3340 10416 3392
rect 10468 3380 10474 3392
rect 10870 3380 10876 3392
rect 10468 3352 10876 3380
rect 10468 3340 10474 3352
rect 10870 3340 10876 3352
rect 10928 3380 10934 3392
rect 11992 3380 12020 3420
rect 12437 3417 12449 3420
rect 12483 3417 12495 3451
rect 12437 3411 12495 3417
rect 10928 3352 12020 3380
rect 13004 3380 13032 3476
rect 13464 3448 13492 3476
rect 14338 3451 14396 3457
rect 14338 3448 14350 3451
rect 13464 3420 14350 3448
rect 14338 3417 14350 3420
rect 14384 3417 14396 3451
rect 16500 3448 16528 3479
rect 16574 3476 16580 3528
rect 16632 3476 16638 3528
rect 16776 3525 16804 3556
rect 16945 3553 16957 3587
rect 16991 3584 17003 3587
rect 18064 3584 18092 3692
rect 18506 3680 18512 3732
rect 18564 3720 18570 3732
rect 18693 3723 18751 3729
rect 18693 3720 18705 3723
rect 18564 3692 18705 3720
rect 18564 3680 18570 3692
rect 18693 3689 18705 3692
rect 18739 3689 18751 3723
rect 18693 3683 18751 3689
rect 20162 3680 20168 3732
rect 20220 3680 20226 3732
rect 18509 3587 18567 3593
rect 18509 3584 18521 3587
rect 16991 3556 18000 3584
rect 18064 3556 18521 3584
rect 16991 3553 17003 3556
rect 16945 3547 17003 3553
rect 16761 3519 16819 3525
rect 16761 3485 16773 3519
rect 16807 3485 16819 3519
rect 16761 3479 16819 3485
rect 17034 3476 17040 3528
rect 17092 3476 17098 3528
rect 17126 3476 17132 3528
rect 17184 3476 17190 3528
rect 17589 3519 17647 3525
rect 17589 3485 17601 3519
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 17681 3519 17739 3525
rect 17681 3485 17693 3519
rect 17727 3516 17739 3519
rect 17770 3516 17776 3528
rect 17727 3488 17776 3516
rect 17727 3485 17739 3488
rect 17681 3479 17739 3485
rect 16666 3448 16672 3460
rect 16500 3420 16672 3448
rect 14338 3411 14396 3417
rect 16666 3408 16672 3420
rect 16724 3448 16730 3460
rect 17052 3448 17080 3476
rect 16724 3420 17080 3448
rect 17604 3448 17632 3479
rect 17770 3476 17776 3488
rect 17828 3476 17834 3528
rect 17972 3525 18000 3556
rect 18509 3553 18521 3556
rect 18555 3553 18567 3587
rect 18509 3547 18567 3553
rect 17957 3519 18015 3525
rect 17957 3485 17969 3519
rect 18003 3485 18015 3519
rect 17957 3479 18015 3485
rect 18138 3476 18144 3528
rect 18196 3516 18202 3528
rect 18877 3519 18935 3525
rect 18877 3516 18889 3519
rect 18196 3488 18889 3516
rect 18196 3476 18202 3488
rect 18877 3485 18889 3488
rect 18923 3485 18935 3519
rect 18877 3479 18935 3485
rect 19061 3519 19119 3525
rect 19061 3485 19073 3519
rect 19107 3516 19119 3519
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 19107 3488 19257 3516
rect 19107 3485 19119 3488
rect 19061 3479 19119 3485
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 19794 3476 19800 3528
rect 19852 3476 19858 3528
rect 19978 3476 19984 3528
rect 20036 3476 20042 3528
rect 17604 3420 17724 3448
rect 16724 3408 16730 3420
rect 13262 3380 13268 3392
rect 13004 3352 13268 3380
rect 10928 3340 10934 3352
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 13446 3340 13452 3392
rect 13504 3340 13510 3392
rect 17696 3380 17724 3420
rect 17862 3408 17868 3460
rect 17920 3448 17926 3460
rect 19812 3448 19840 3476
rect 17920 3420 19840 3448
rect 17920 3408 17926 3420
rect 18046 3380 18052 3392
rect 17696 3352 18052 3380
rect 18046 3340 18052 3352
rect 18104 3380 18110 3392
rect 18506 3380 18512 3392
rect 18104 3352 18512 3380
rect 18104 3340 18110 3352
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 1104 3290 22264 3312
rect 1104 3238 4255 3290
rect 4307 3238 4319 3290
rect 4371 3238 4383 3290
rect 4435 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 9545 3290
rect 9597 3238 9609 3290
rect 9661 3238 9673 3290
rect 9725 3238 9737 3290
rect 9789 3238 9801 3290
rect 9853 3238 14835 3290
rect 14887 3238 14899 3290
rect 14951 3238 14963 3290
rect 15015 3238 15027 3290
rect 15079 3238 15091 3290
rect 15143 3238 20125 3290
rect 20177 3238 20189 3290
rect 20241 3238 20253 3290
rect 20305 3238 20317 3290
rect 20369 3238 20381 3290
rect 20433 3238 22264 3290
rect 1104 3216 22264 3238
rect 4614 3136 4620 3188
rect 4672 3136 4678 3188
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 5997 3179 6055 3185
rect 5997 3176 6009 3179
rect 5224 3148 6009 3176
rect 5224 3136 5230 3148
rect 5997 3145 6009 3148
rect 6043 3145 6055 3179
rect 5997 3139 6055 3145
rect 6086 3136 6092 3188
rect 6144 3136 6150 3188
rect 6270 3136 6276 3188
rect 6328 3176 6334 3188
rect 6523 3179 6581 3185
rect 6523 3176 6535 3179
rect 6328 3148 6535 3176
rect 6328 3136 6334 3148
rect 6523 3145 6535 3148
rect 6569 3145 6581 3179
rect 6822 3176 6828 3188
rect 6523 3139 6581 3145
rect 6656 3148 6828 3176
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4212 3012 4445 3040
rect 4212 3000 4218 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4632 3040 4660 3136
rect 6104 3108 6132 3136
rect 5920 3080 6132 3108
rect 5920 3049 5948 3080
rect 4689 3043 4747 3049
rect 4689 3040 4701 3043
rect 4632 3012 4701 3040
rect 4433 3003 4491 3009
rect 4689 3009 4701 3012
rect 4735 3009 4747 3043
rect 4689 3003 4747 3009
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 6089 3043 6147 3049
rect 6089 3009 6101 3043
rect 6135 3040 6147 3043
rect 6656 3040 6684 3148
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 8202 3176 8208 3188
rect 8128 3148 8208 3176
rect 6733 3111 6791 3117
rect 6733 3077 6745 3111
rect 6779 3108 6791 3111
rect 6932 3108 6960 3136
rect 6779 3080 6960 3108
rect 7960 3111 8018 3117
rect 6779 3077 6791 3080
rect 6733 3071 6791 3077
rect 7960 3077 7972 3111
rect 8006 3108 8018 3111
rect 8128 3108 8156 3148
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8294 3136 8300 3188
rect 8352 3136 8358 3188
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 8435 3148 9168 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 8312 3108 8340 3136
rect 8006 3080 8156 3108
rect 8220 3080 8984 3108
rect 8006 3077 8018 3080
rect 7960 3071 8018 3077
rect 8220 3049 8248 3080
rect 8205 3043 8263 3049
rect 6135 3012 6500 3040
rect 6656 3012 8156 3040
rect 6135 3009 6147 3012
rect 6089 3003 6147 3009
rect 5813 2907 5871 2913
rect 5813 2873 5825 2907
rect 5859 2904 5871 2907
rect 5902 2904 5908 2916
rect 5859 2876 5908 2904
rect 5859 2873 5871 2876
rect 5813 2867 5871 2873
rect 5902 2864 5908 2876
rect 5960 2904 5966 2916
rect 6270 2904 6276 2916
rect 5960 2876 6276 2904
rect 5960 2864 5966 2876
rect 6270 2864 6276 2876
rect 6328 2864 6334 2916
rect 6472 2904 6500 3012
rect 8128 2972 8156 3012
rect 8205 3009 8217 3043
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 8312 2972 8340 3003
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 8956 3049 8984 3080
rect 8573 3043 8631 3049
rect 8573 3040 8585 3043
rect 8536 3012 8585 3040
rect 8536 3000 8542 3012
rect 8573 3009 8585 3012
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3009 8999 3043
rect 9140 3040 9168 3148
rect 10042 3136 10048 3188
rect 10100 3136 10106 3188
rect 10321 3179 10379 3185
rect 10321 3145 10333 3179
rect 10367 3176 10379 3179
rect 11146 3176 11152 3188
rect 10367 3148 11152 3176
rect 10367 3145 10379 3148
rect 10321 3139 10379 3145
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 11517 3179 11575 3185
rect 11517 3145 11529 3179
rect 11563 3176 11575 3179
rect 12434 3176 12440 3188
rect 11563 3148 12440 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 9208 3111 9266 3117
rect 9208 3077 9220 3111
rect 9254 3108 9266 3111
rect 10060 3108 10088 3136
rect 9254 3080 10088 3108
rect 9254 3077 9266 3080
rect 9208 3071 9266 3077
rect 10778 3068 10784 3120
rect 10836 3068 10842 3120
rect 9490 3040 9496 3052
rect 9140 3012 9496 3040
rect 8941 3003 8999 3009
rect 9490 3000 9496 3012
rect 9548 3040 9554 3052
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 9548 3012 10517 3040
rect 9548 3000 9554 3012
rect 10505 3009 10517 3012
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3040 10655 3043
rect 10796 3040 10824 3068
rect 11054 3049 11060 3052
rect 10643 3012 10824 3040
rect 11035 3043 11060 3049
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 11035 3009 11047 3043
rect 11035 3003 11060 3009
rect 11054 3000 11060 3003
rect 11112 3000 11118 3052
rect 11238 3000 11244 3052
rect 11296 3000 11302 3052
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3040 11391 3043
rect 11532 3040 11560 3139
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 14277 3179 14335 3185
rect 14277 3145 14289 3179
rect 14323 3176 14335 3179
rect 14734 3176 14740 3188
rect 14323 3148 14740 3176
rect 14323 3145 14335 3148
rect 14277 3139 14335 3145
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 16117 3179 16175 3185
rect 16117 3145 16129 3179
rect 16163 3145 16175 3179
rect 16117 3139 16175 3145
rect 11790 3068 11796 3120
rect 11848 3068 11854 3120
rect 12066 3068 12072 3120
rect 12124 3108 12130 3120
rect 12345 3111 12403 3117
rect 12345 3108 12357 3111
rect 12124 3080 12357 3108
rect 12124 3068 12130 3080
rect 12345 3077 12357 3080
rect 12391 3077 12403 3111
rect 12345 3071 12403 3077
rect 11379 3012 11560 3040
rect 11379 3009 11391 3012
rect 11333 3003 11391 3009
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11664 3012 11713 3040
rect 11664 3000 11670 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11808 3040 11836 3068
rect 12452 3049 12480 3136
rect 14912 3111 14970 3117
rect 12912 3080 14688 3108
rect 12912 3052 12940 3080
rect 11885 3043 11943 3049
rect 11885 3040 11897 3043
rect 11808 3012 11897 3040
rect 11701 3003 11759 3009
rect 11885 3009 11897 3012
rect 11931 3040 11943 3043
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11931 3012 11989 3040
rect 11931 3009 11943 3012
rect 11885 3003 11943 3009
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3009 12219 3043
rect 12161 3003 12219 3009
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3009 12495 3043
rect 12437 3003 12495 3009
rect 11149 2975 11207 2981
rect 8128 2944 8340 2972
rect 10612 2944 11100 2972
rect 10612 2916 10640 2944
rect 6472 2876 7328 2904
rect 6365 2839 6423 2845
rect 6365 2805 6377 2839
rect 6411 2836 6423 2839
rect 6472 2836 6500 2876
rect 6411 2808 6500 2836
rect 6411 2805 6423 2808
rect 6365 2799 6423 2805
rect 6546 2796 6552 2848
rect 6604 2796 6610 2848
rect 7300 2836 7328 2876
rect 10594 2864 10600 2916
rect 10652 2864 10658 2916
rect 10870 2864 10876 2916
rect 10928 2904 10934 2916
rect 10965 2907 11023 2913
rect 10965 2904 10977 2907
rect 10928 2876 10977 2904
rect 10928 2864 10934 2876
rect 10965 2873 10977 2876
rect 11011 2873 11023 2907
rect 11072 2904 11100 2944
rect 11149 2941 11161 2975
rect 11195 2972 11207 2975
rect 11256 2972 11284 3000
rect 11716 2972 11744 3003
rect 12176 2972 12204 3003
rect 12894 3000 12900 3052
rect 12952 3000 12958 3052
rect 13170 3049 13176 3052
rect 13164 3003 13176 3049
rect 13170 3000 13176 3003
rect 13228 3000 13234 3052
rect 14660 3049 14688 3080
rect 14912 3077 14924 3111
rect 14958 3108 14970 3111
rect 16132 3108 16160 3139
rect 16206 3136 16212 3188
rect 16264 3136 16270 3188
rect 16390 3136 16396 3188
rect 16448 3176 16454 3188
rect 16669 3179 16727 3185
rect 16669 3176 16681 3179
rect 16448 3148 16681 3176
rect 16448 3136 16454 3148
rect 16669 3145 16681 3148
rect 16715 3145 16727 3179
rect 16669 3139 16727 3145
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 18138 3176 18144 3188
rect 17184 3148 18144 3176
rect 17184 3136 17190 3148
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 19334 3136 19340 3188
rect 19392 3136 19398 3188
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 20349 3179 20407 3185
rect 20349 3176 20361 3179
rect 20036 3148 20361 3176
rect 20036 3136 20042 3148
rect 20349 3145 20361 3148
rect 20395 3145 20407 3179
rect 20349 3139 20407 3145
rect 14958 3080 16160 3108
rect 14958 3077 14970 3080
rect 14912 3071 14970 3077
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3009 14703 3043
rect 16224 3040 16252 3136
rect 19352 3108 19380 3136
rect 18064 3080 19564 3108
rect 16301 3043 16359 3049
rect 16301 3040 16313 3043
rect 16224 3012 16313 3040
rect 14645 3003 14703 3009
rect 16301 3009 16313 3012
rect 16347 3009 16359 3043
rect 16301 3003 16359 3009
rect 17494 3000 17500 3052
rect 17552 3040 17558 3052
rect 18064 3049 18092 3080
rect 17782 3043 17840 3049
rect 17782 3040 17794 3043
rect 17552 3012 17794 3040
rect 17552 3000 17558 3012
rect 17782 3009 17794 3012
rect 17828 3009 17840 3043
rect 17782 3003 17840 3009
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 18874 3000 18880 3052
rect 18932 3040 18938 3052
rect 19536 3049 19564 3080
rect 19254 3043 19312 3049
rect 19254 3040 19266 3043
rect 18932 3012 19266 3040
rect 18932 3000 18938 3012
rect 19254 3009 19266 3012
rect 19300 3009 19312 3043
rect 19254 3003 19312 3009
rect 19521 3043 19579 3049
rect 19521 3009 19533 3043
rect 19567 3009 19579 3043
rect 19521 3003 19579 3009
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3040 20223 3043
rect 21450 3040 21456 3052
rect 20211 3012 21456 3040
rect 20211 3009 20223 3012
rect 20165 3003 20223 3009
rect 21450 3000 21456 3012
rect 21508 3000 21514 3052
rect 11195 2944 11284 2972
rect 11440 2944 11652 2972
rect 11716 2944 12204 2972
rect 11195 2941 11207 2944
rect 11149 2935 11207 2941
rect 11241 2907 11299 2913
rect 11241 2904 11253 2907
rect 11072 2876 11253 2904
rect 10965 2867 11023 2873
rect 11241 2873 11253 2876
rect 11287 2904 11299 2907
rect 11440 2904 11468 2944
rect 11287 2876 11468 2904
rect 11624 2904 11652 2944
rect 16666 2932 16672 2984
rect 16724 2932 16730 2984
rect 19981 2975 20039 2981
rect 19981 2941 19993 2975
rect 20027 2941 20039 2975
rect 19981 2935 20039 2941
rect 12158 2904 12164 2916
rect 11624 2876 12164 2904
rect 11287 2873 11299 2876
rect 11241 2867 11299 2873
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 16025 2907 16083 2913
rect 16025 2873 16037 2907
rect 16071 2904 16083 2907
rect 16684 2904 16712 2932
rect 16071 2876 16712 2904
rect 18064 2876 18644 2904
rect 16071 2873 16083 2876
rect 16025 2867 16083 2873
rect 8018 2836 8024 2848
rect 7300 2808 8024 2836
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 8570 2796 8576 2848
rect 8628 2796 8634 2848
rect 9214 2796 9220 2848
rect 9272 2836 9278 2848
rect 11606 2836 11612 2848
rect 9272 2808 11612 2836
rect 9272 2796 9278 2808
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 18064 2836 18092 2876
rect 13320 2808 18092 2836
rect 18141 2839 18199 2845
rect 13320 2796 13326 2808
rect 18141 2805 18153 2839
rect 18187 2836 18199 2839
rect 18506 2836 18512 2848
rect 18187 2808 18512 2836
rect 18187 2805 18199 2808
rect 18141 2799 18199 2805
rect 18506 2796 18512 2808
rect 18564 2796 18570 2848
rect 18616 2836 18644 2876
rect 19996 2836 20024 2935
rect 18616 2808 20024 2836
rect 1104 2746 22264 2768
rect 1104 2694 3595 2746
rect 3647 2694 3659 2746
rect 3711 2694 3723 2746
rect 3775 2694 3787 2746
rect 3839 2694 3851 2746
rect 3903 2694 8885 2746
rect 8937 2694 8949 2746
rect 9001 2694 9013 2746
rect 9065 2694 9077 2746
rect 9129 2694 9141 2746
rect 9193 2694 14175 2746
rect 14227 2694 14239 2746
rect 14291 2694 14303 2746
rect 14355 2694 14367 2746
rect 14419 2694 14431 2746
rect 14483 2694 19465 2746
rect 19517 2694 19529 2746
rect 19581 2694 19593 2746
rect 19645 2694 19657 2746
rect 19709 2694 19721 2746
rect 19773 2694 22264 2746
rect 1104 2672 22264 2694
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 13357 2635 13415 2641
rect 13357 2632 13369 2635
rect 13228 2604 13369 2632
rect 13228 2592 13234 2604
rect 13357 2601 13369 2604
rect 13403 2601 13415 2635
rect 13357 2595 13415 2601
rect 17129 2635 17187 2641
rect 17129 2601 17141 2635
rect 17175 2632 17187 2635
rect 17494 2632 17500 2644
rect 17175 2604 17500 2632
rect 17175 2601 17187 2604
rect 17129 2595 17187 2601
rect 17494 2592 17500 2604
rect 17552 2592 17558 2644
rect 17954 2592 17960 2644
rect 18012 2592 18018 2644
rect 18874 2592 18880 2644
rect 18932 2592 18938 2644
rect 18966 2592 18972 2644
rect 19024 2632 19030 2644
rect 19245 2635 19303 2641
rect 19245 2632 19257 2635
rect 19024 2604 19257 2632
rect 19024 2592 19030 2604
rect 19245 2601 19257 2604
rect 19291 2601 19303 2635
rect 19245 2595 19303 2601
rect 21450 2592 21456 2644
rect 21508 2592 21514 2644
rect 17972 2564 18000 2592
rect 17972 2536 18736 2564
rect 17126 2456 17132 2508
rect 17184 2496 17190 2508
rect 17184 2468 17632 2496
rect 17184 2456 17190 2468
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 9033 2431 9091 2437
rect 9033 2428 9045 2431
rect 8628 2400 9045 2428
rect 8628 2388 8634 2400
rect 9033 2397 9045 2400
rect 9079 2397 9091 2431
rect 9033 2391 9091 2397
rect 13538 2388 13544 2440
rect 13596 2388 13602 2440
rect 17604 2437 17632 2468
rect 18506 2456 18512 2508
rect 18564 2456 18570 2508
rect 18708 2437 18736 2536
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2428 17003 2431
rect 17405 2431 17463 2437
rect 17405 2428 17417 2431
rect 16991 2400 17417 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 17405 2397 17417 2400
rect 17451 2397 17463 2431
rect 17405 2391 17463 2397
rect 17589 2431 17647 2437
rect 17589 2397 17601 2431
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2428 17831 2431
rect 17957 2431 18015 2437
rect 17957 2428 17969 2431
rect 17819 2400 17969 2428
rect 17819 2397 17831 2400
rect 17773 2391 17831 2397
rect 17957 2397 17969 2400
rect 18003 2397 18015 2431
rect 17957 2391 18015 2397
rect 18693 2431 18751 2437
rect 18693 2397 18705 2431
rect 18739 2397 18751 2431
rect 18693 2391 18751 2397
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 21637 2431 21695 2437
rect 21637 2397 21649 2431
rect 21683 2428 21695 2431
rect 21683 2400 22232 2428
rect 21683 2397 21695 2400
rect 21637 2391 21695 2397
rect 6886 2332 13124 2360
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2292 1639 2295
rect 6886 2292 6914 2332
rect 13096 2304 13124 2332
rect 17862 2320 17868 2372
rect 17920 2360 17926 2372
rect 19444 2360 19472 2391
rect 17920 2332 19472 2360
rect 17920 2320 17926 2332
rect 22204 2304 22232 2400
rect 1627 2264 6914 2292
rect 1627 2261 1639 2264
rect 1581 2255 1639 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8444 2264 9137 2292
rect 8444 2252 8450 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 13078 2252 13084 2304
rect 13136 2252 13142 2304
rect 22186 2252 22192 2304
rect 22244 2252 22250 2304
rect 1104 2202 22264 2224
rect 1104 2150 4255 2202
rect 4307 2150 4319 2202
rect 4371 2150 4383 2202
rect 4435 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 9545 2202
rect 9597 2150 9609 2202
rect 9661 2150 9673 2202
rect 9725 2150 9737 2202
rect 9789 2150 9801 2202
rect 9853 2150 14835 2202
rect 14887 2150 14899 2202
rect 14951 2150 14963 2202
rect 15015 2150 15027 2202
rect 15079 2150 15091 2202
rect 15143 2150 20125 2202
rect 20177 2150 20189 2202
rect 20241 2150 20253 2202
rect 20305 2150 20317 2202
rect 20369 2150 20381 2202
rect 20433 2150 22264 2202
rect 1104 2128 22264 2150
<< via1 >>
rect 4255 22822 4307 22874
rect 4319 22822 4371 22874
rect 4383 22822 4435 22874
rect 4447 22822 4499 22874
rect 4511 22822 4563 22874
rect 9545 22822 9597 22874
rect 9609 22822 9661 22874
rect 9673 22822 9725 22874
rect 9737 22822 9789 22874
rect 9801 22822 9853 22874
rect 14835 22822 14887 22874
rect 14899 22822 14951 22874
rect 14963 22822 15015 22874
rect 15027 22822 15079 22874
rect 15091 22822 15143 22874
rect 20125 22822 20177 22874
rect 20189 22822 20241 22874
rect 20253 22822 20305 22874
rect 20317 22822 20369 22874
rect 20381 22822 20433 22874
rect 1308 22720 1360 22772
rect 10324 22720 10376 22772
rect 19340 22720 19392 22772
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 13452 22627 13504 22636
rect 13452 22593 13461 22627
rect 13461 22593 13495 22627
rect 13495 22593 13504 22627
rect 13452 22584 13504 22593
rect 13636 22627 13688 22636
rect 13636 22593 13645 22627
rect 13645 22593 13679 22627
rect 13679 22593 13688 22627
rect 13636 22584 13688 22593
rect 13544 22516 13596 22568
rect 16764 22627 16816 22636
rect 16764 22593 16773 22627
rect 16773 22593 16807 22627
rect 16807 22593 16816 22627
rect 16764 22584 16816 22593
rect 16948 22423 17000 22432
rect 16948 22389 16957 22423
rect 16957 22389 16991 22423
rect 16991 22389 17000 22423
rect 16948 22380 17000 22389
rect 19340 22380 19392 22432
rect 3595 22278 3647 22330
rect 3659 22278 3711 22330
rect 3723 22278 3775 22330
rect 3787 22278 3839 22330
rect 3851 22278 3903 22330
rect 8885 22278 8937 22330
rect 8949 22278 9001 22330
rect 9013 22278 9065 22330
rect 9077 22278 9129 22330
rect 9141 22278 9193 22330
rect 14175 22278 14227 22330
rect 14239 22278 14291 22330
rect 14303 22278 14355 22330
rect 14367 22278 14419 22330
rect 14431 22278 14483 22330
rect 19465 22278 19517 22330
rect 19529 22278 19581 22330
rect 19593 22278 19645 22330
rect 19657 22278 19709 22330
rect 19721 22278 19773 22330
rect 7564 22108 7616 22160
rect 8392 22108 8444 22160
rect 12992 22108 13044 22160
rect 2596 22040 2648 22092
rect 4896 22040 4948 22092
rect 3424 21972 3476 22024
rect 2964 21947 3016 21956
rect 2964 21913 2973 21947
rect 2973 21913 3007 21947
rect 3007 21913 3016 21947
rect 2964 21904 3016 21913
rect 6736 21972 6788 22024
rect 5724 21904 5776 21956
rect 7380 21904 7432 21956
rect 3056 21879 3108 21888
rect 3056 21845 3071 21879
rect 3071 21845 3105 21879
rect 3105 21845 3108 21879
rect 3056 21836 3108 21845
rect 3516 21836 3568 21888
rect 4068 21836 4120 21888
rect 7104 21836 7156 21888
rect 7196 21836 7248 21888
rect 8300 22015 8352 22024
rect 8300 21981 8309 22015
rect 8309 21981 8343 22015
rect 8343 21981 8352 22015
rect 8300 21972 8352 21981
rect 9956 22015 10008 22024
rect 9956 21981 9965 22015
rect 9965 21981 9999 22015
rect 9999 21981 10008 22015
rect 9956 21972 10008 21981
rect 12716 22040 12768 22092
rect 10416 21904 10468 21956
rect 7748 21836 7800 21888
rect 7840 21879 7892 21888
rect 7840 21845 7849 21879
rect 7849 21845 7883 21879
rect 7883 21845 7892 21879
rect 7840 21836 7892 21845
rect 8484 21879 8536 21888
rect 8484 21845 8493 21879
rect 8493 21845 8527 21879
rect 8527 21845 8536 21879
rect 8484 21836 8536 21845
rect 12072 21972 12124 22024
rect 13084 22015 13136 22024
rect 13084 21981 13093 22015
rect 13093 21981 13127 22015
rect 13127 21981 13136 22015
rect 13084 21972 13136 21981
rect 12164 21947 12216 21956
rect 12164 21913 12173 21947
rect 12173 21913 12207 21947
rect 12207 21913 12216 21947
rect 12164 21904 12216 21913
rect 12348 21947 12400 21956
rect 12348 21913 12357 21947
rect 12357 21913 12391 21947
rect 12391 21913 12400 21947
rect 12348 21904 12400 21913
rect 11428 21879 11480 21888
rect 11428 21845 11437 21879
rect 11437 21845 11471 21879
rect 11471 21845 11480 21879
rect 11428 21836 11480 21845
rect 12072 21836 12124 21888
rect 13636 21836 13688 21888
rect 13728 21879 13780 21888
rect 13728 21845 13737 21879
rect 13737 21845 13771 21879
rect 13771 21845 13780 21879
rect 13728 21836 13780 21845
rect 14280 21904 14332 21956
rect 19064 21972 19116 22024
rect 16948 21904 17000 21956
rect 15292 21836 15344 21888
rect 4255 21734 4307 21786
rect 4319 21734 4371 21786
rect 4383 21734 4435 21786
rect 4447 21734 4499 21786
rect 4511 21734 4563 21786
rect 9545 21734 9597 21786
rect 9609 21734 9661 21786
rect 9673 21734 9725 21786
rect 9737 21734 9789 21786
rect 9801 21734 9853 21786
rect 14835 21734 14887 21786
rect 14899 21734 14951 21786
rect 14963 21734 15015 21786
rect 15027 21734 15079 21786
rect 15091 21734 15143 21786
rect 20125 21734 20177 21786
rect 20189 21734 20241 21786
rect 20253 21734 20305 21786
rect 20317 21734 20369 21786
rect 20381 21734 20433 21786
rect 1768 21428 1820 21480
rect 2504 21539 2556 21548
rect 2504 21505 2513 21539
rect 2513 21505 2547 21539
rect 2547 21505 2556 21539
rect 2504 21496 2556 21505
rect 3056 21632 3108 21684
rect 5724 21675 5776 21684
rect 5724 21641 5733 21675
rect 5733 21641 5767 21675
rect 5767 21641 5776 21675
rect 5724 21632 5776 21641
rect 6828 21632 6880 21684
rect 7196 21632 7248 21684
rect 10416 21675 10468 21684
rect 10416 21641 10425 21675
rect 10425 21641 10459 21675
rect 10459 21641 10468 21675
rect 10416 21632 10468 21641
rect 11428 21632 11480 21684
rect 11888 21632 11940 21684
rect 12072 21632 12124 21684
rect 13084 21675 13136 21684
rect 13084 21641 13093 21675
rect 13093 21641 13127 21675
rect 13127 21641 13136 21675
rect 13084 21632 13136 21641
rect 13452 21632 13504 21684
rect 13728 21632 13780 21684
rect 14280 21675 14332 21684
rect 14280 21641 14289 21675
rect 14289 21641 14323 21675
rect 14323 21641 14332 21675
rect 14280 21632 14332 21641
rect 6092 21607 6144 21616
rect 6092 21573 6101 21607
rect 6101 21573 6135 21607
rect 6135 21573 6144 21607
rect 6092 21564 6144 21573
rect 2596 21360 2648 21412
rect 4068 21403 4120 21412
rect 4068 21369 4077 21403
rect 4077 21369 4111 21403
rect 4111 21369 4120 21403
rect 4068 21360 4120 21369
rect 6184 21539 6236 21548
rect 6184 21505 6193 21539
rect 6193 21505 6227 21539
rect 6227 21505 6236 21539
rect 6184 21496 6236 21505
rect 6736 21496 6788 21548
rect 7840 21564 7892 21616
rect 8484 21564 8536 21616
rect 7104 21496 7156 21548
rect 6276 21428 6328 21480
rect 6920 21428 6972 21480
rect 7564 21428 7616 21480
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 13452 21539 13504 21548
rect 13452 21505 13461 21539
rect 13461 21505 13495 21539
rect 13495 21505 13504 21539
rect 13452 21496 13504 21505
rect 13636 21496 13688 21548
rect 15292 21564 15344 21616
rect 5724 21360 5776 21412
rect 3976 21292 4028 21344
rect 5540 21292 5592 21344
rect 6644 21292 6696 21344
rect 6736 21335 6788 21344
rect 6736 21301 6745 21335
rect 6745 21301 6779 21335
rect 6779 21301 6788 21335
rect 6736 21292 6788 21301
rect 7104 21335 7156 21344
rect 7104 21301 7113 21335
rect 7113 21301 7147 21335
rect 7147 21301 7156 21335
rect 7104 21292 7156 21301
rect 13544 21428 13596 21480
rect 14004 21471 14056 21480
rect 14004 21437 14013 21471
rect 14013 21437 14047 21471
rect 14047 21437 14056 21471
rect 14004 21428 14056 21437
rect 14096 21471 14148 21480
rect 14096 21437 14105 21471
rect 14105 21437 14139 21471
rect 14139 21437 14148 21471
rect 14096 21428 14148 21437
rect 16580 21632 16632 21684
rect 15844 21539 15896 21548
rect 15844 21505 15853 21539
rect 15853 21505 15887 21539
rect 15887 21505 15896 21539
rect 15844 21496 15896 21505
rect 16028 21539 16080 21548
rect 16028 21505 16037 21539
rect 16037 21505 16071 21539
rect 16071 21505 16080 21539
rect 16028 21496 16080 21505
rect 16120 21539 16172 21548
rect 16120 21505 16129 21539
rect 16129 21505 16163 21539
rect 16163 21505 16172 21539
rect 16120 21496 16172 21505
rect 15200 21428 15252 21480
rect 15292 21428 15344 21480
rect 16672 21539 16724 21548
rect 16672 21505 16681 21539
rect 16681 21505 16715 21539
rect 16715 21505 16724 21539
rect 16672 21496 16724 21505
rect 22192 21496 22244 21548
rect 15016 21360 15068 21412
rect 16948 21360 17000 21412
rect 9864 21292 9916 21344
rect 10784 21335 10836 21344
rect 10784 21301 10793 21335
rect 10793 21301 10827 21335
rect 10827 21301 10836 21335
rect 10784 21292 10836 21301
rect 14924 21335 14976 21344
rect 14924 21301 14933 21335
rect 14933 21301 14967 21335
rect 14967 21301 14976 21335
rect 14924 21292 14976 21301
rect 15476 21292 15528 21344
rect 16304 21335 16356 21344
rect 16304 21301 16313 21335
rect 16313 21301 16347 21335
rect 16347 21301 16356 21335
rect 16304 21292 16356 21301
rect 16764 21335 16816 21344
rect 16764 21301 16773 21335
rect 16773 21301 16807 21335
rect 16807 21301 16816 21335
rect 16764 21292 16816 21301
rect 16856 21292 16908 21344
rect 20628 21292 20680 21344
rect 3595 21190 3647 21242
rect 3659 21190 3711 21242
rect 3723 21190 3775 21242
rect 3787 21190 3839 21242
rect 3851 21190 3903 21242
rect 8885 21190 8937 21242
rect 8949 21190 9001 21242
rect 9013 21190 9065 21242
rect 9077 21190 9129 21242
rect 9141 21190 9193 21242
rect 14175 21190 14227 21242
rect 14239 21190 14291 21242
rect 14303 21190 14355 21242
rect 14367 21190 14419 21242
rect 14431 21190 14483 21242
rect 19465 21190 19517 21242
rect 19529 21190 19581 21242
rect 19593 21190 19645 21242
rect 19657 21190 19709 21242
rect 19721 21190 19773 21242
rect 2504 21088 2556 21140
rect 2964 21088 3016 21140
rect 3424 21131 3476 21140
rect 3424 21097 3433 21131
rect 3433 21097 3467 21131
rect 3467 21097 3476 21131
rect 3424 21088 3476 21097
rect 3516 21088 3568 21140
rect 3976 21088 4028 21140
rect 4068 21088 4120 21140
rect 6184 21088 6236 21140
rect 6276 21088 6328 21140
rect 6736 21088 6788 21140
rect 6828 21088 6880 21140
rect 7380 21088 7432 21140
rect 7748 21131 7800 21140
rect 7748 21097 7757 21131
rect 7757 21097 7791 21131
rect 7791 21097 7800 21131
rect 7748 21088 7800 21097
rect 7840 21088 7892 21140
rect 8300 21131 8352 21140
rect 8300 21097 8309 21131
rect 8309 21097 8343 21131
rect 8343 21097 8352 21131
rect 8300 21088 8352 21097
rect 8484 21131 8536 21140
rect 8484 21097 8493 21131
rect 8493 21097 8527 21131
rect 8527 21097 8536 21131
rect 8484 21088 8536 21097
rect 10416 21088 10468 21140
rect 11980 21131 12032 21140
rect 11980 21097 11989 21131
rect 11989 21097 12023 21131
rect 12023 21097 12032 21131
rect 11980 21088 12032 21097
rect 3148 20884 3200 20936
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 4068 20927 4120 20936
rect 4068 20893 4077 20927
rect 4077 20893 4111 20927
rect 4111 20893 4120 20927
rect 4068 20884 4120 20893
rect 5540 20952 5592 21004
rect 6092 20952 6144 21004
rect 5816 20884 5868 20936
rect 5908 20927 5960 20936
rect 5908 20893 5917 20927
rect 5917 20893 5951 20927
rect 5951 20893 5960 20927
rect 5908 20884 5960 20893
rect 6644 20995 6696 21004
rect 6644 20961 6653 20995
rect 6653 20961 6687 20995
rect 6687 20961 6696 20995
rect 6644 20952 6696 20961
rect 5816 20748 5868 20800
rect 6828 20748 6880 20800
rect 12256 21088 12308 21140
rect 12716 21088 12768 21140
rect 12992 21131 13044 21140
rect 12992 21097 13001 21131
rect 13001 21097 13035 21131
rect 13035 21097 13044 21131
rect 12992 21088 13044 21097
rect 13084 21088 13136 21140
rect 13544 21088 13596 21140
rect 14096 21088 14148 21140
rect 14924 21088 14976 21140
rect 15016 21088 15068 21140
rect 15476 21088 15528 21140
rect 7564 20927 7616 20936
rect 7564 20893 7573 20927
rect 7573 20893 7607 20927
rect 7607 20893 7616 20927
rect 7564 20884 7616 20893
rect 7656 20927 7708 20936
rect 7656 20893 7665 20927
rect 7665 20893 7699 20927
rect 7699 20893 7708 20927
rect 7656 20884 7708 20893
rect 7748 20859 7800 20868
rect 7748 20825 7757 20859
rect 7757 20825 7791 20859
rect 7791 20825 7800 20859
rect 7748 20816 7800 20825
rect 8668 20859 8720 20868
rect 8668 20825 8677 20859
rect 8677 20825 8711 20859
rect 8711 20825 8720 20859
rect 8668 20816 8720 20825
rect 9312 20748 9364 20800
rect 9864 20884 9916 20936
rect 10784 20884 10836 20936
rect 10232 20816 10284 20868
rect 15568 21020 15620 21072
rect 15844 21088 15896 21140
rect 16120 21088 16172 21140
rect 16396 21088 16448 21140
rect 16764 21088 16816 21140
rect 15752 20995 15804 21004
rect 15752 20961 15761 20995
rect 15761 20961 15795 20995
rect 15795 20961 15804 20995
rect 15752 20952 15804 20961
rect 16028 21020 16080 21072
rect 15568 20927 15620 20936
rect 15568 20893 15577 20927
rect 15577 20893 15611 20927
rect 15611 20893 15620 20927
rect 15568 20884 15620 20893
rect 10324 20748 10376 20800
rect 10968 20748 11020 20800
rect 11152 20748 11204 20800
rect 11244 20791 11296 20800
rect 11244 20757 11253 20791
rect 11253 20757 11287 20791
rect 11287 20757 11296 20791
rect 11244 20748 11296 20757
rect 13084 20748 13136 20800
rect 15476 20748 15528 20800
rect 15752 20748 15804 20800
rect 4255 20646 4307 20698
rect 4319 20646 4371 20698
rect 4383 20646 4435 20698
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 9545 20646 9597 20698
rect 9609 20646 9661 20698
rect 9673 20646 9725 20698
rect 9737 20646 9789 20698
rect 9801 20646 9853 20698
rect 14835 20646 14887 20698
rect 14899 20646 14951 20698
rect 14963 20646 15015 20698
rect 15027 20646 15079 20698
rect 15091 20646 15143 20698
rect 20125 20646 20177 20698
rect 20189 20646 20241 20698
rect 20253 20646 20305 20698
rect 20317 20646 20369 20698
rect 20381 20646 20433 20698
rect 3976 20544 4028 20596
rect 5908 20544 5960 20596
rect 6920 20544 6972 20596
rect 7104 20544 7156 20596
rect 7288 20544 7340 20596
rect 7748 20544 7800 20596
rect 10232 20587 10284 20596
rect 10232 20553 10241 20587
rect 10241 20553 10275 20587
rect 10275 20553 10284 20587
rect 10232 20544 10284 20553
rect 10784 20587 10836 20596
rect 10784 20553 10793 20587
rect 10793 20553 10827 20587
rect 10827 20553 10836 20587
rect 10784 20544 10836 20553
rect 12164 20544 12216 20596
rect 12256 20544 12308 20596
rect 8668 20476 8720 20528
rect 11336 20476 11388 20528
rect 15292 20587 15344 20596
rect 15292 20553 15301 20587
rect 15301 20553 15335 20587
rect 15335 20553 15344 20587
rect 15292 20544 15344 20553
rect 15568 20544 15620 20596
rect 6736 20451 6788 20460
rect 6736 20417 6745 20451
rect 6745 20417 6779 20451
rect 6779 20417 6788 20451
rect 6736 20408 6788 20417
rect 6828 20408 6880 20460
rect 10416 20451 10468 20460
rect 10416 20417 10425 20451
rect 10425 20417 10459 20451
rect 10459 20417 10468 20451
rect 10416 20408 10468 20417
rect 10968 20451 11020 20460
rect 10968 20417 10977 20451
rect 10977 20417 11011 20451
rect 11011 20417 11020 20451
rect 10968 20408 11020 20417
rect 11244 20408 11296 20460
rect 12072 20408 12124 20460
rect 12348 20408 12400 20460
rect 15200 20451 15252 20460
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 15752 20451 15804 20460
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 3976 20272 4028 20324
rect 16212 20340 16264 20392
rect 16396 20451 16448 20460
rect 16396 20417 16405 20451
rect 16405 20417 16439 20451
rect 16439 20417 16448 20451
rect 16396 20408 16448 20417
rect 20628 20544 20680 20596
rect 16948 20451 17000 20460
rect 16948 20417 16957 20451
rect 16957 20417 16991 20451
rect 16991 20417 17000 20451
rect 16948 20408 17000 20417
rect 3148 20204 3200 20256
rect 12256 20272 12308 20324
rect 16672 20315 16724 20324
rect 16672 20281 16681 20315
rect 16681 20281 16715 20315
rect 16715 20281 16724 20315
rect 16672 20272 16724 20281
rect 11152 20204 11204 20256
rect 12532 20247 12584 20256
rect 12532 20213 12541 20247
rect 12541 20213 12575 20247
rect 12575 20213 12584 20247
rect 12532 20204 12584 20213
rect 15476 20204 15528 20256
rect 16120 20204 16172 20256
rect 16396 20204 16448 20256
rect 20168 20204 20220 20256
rect 20536 20247 20588 20256
rect 20536 20213 20545 20247
rect 20545 20213 20579 20247
rect 20579 20213 20588 20247
rect 20536 20204 20588 20213
rect 3595 20102 3647 20154
rect 3659 20102 3711 20154
rect 3723 20102 3775 20154
rect 3787 20102 3839 20154
rect 3851 20102 3903 20154
rect 8885 20102 8937 20154
rect 8949 20102 9001 20154
rect 9013 20102 9065 20154
rect 9077 20102 9129 20154
rect 9141 20102 9193 20154
rect 14175 20102 14227 20154
rect 14239 20102 14291 20154
rect 14303 20102 14355 20154
rect 14367 20102 14419 20154
rect 14431 20102 14483 20154
rect 19465 20102 19517 20154
rect 19529 20102 19581 20154
rect 19593 20102 19645 20154
rect 19657 20102 19709 20154
rect 19721 20102 19773 20154
rect 3240 19796 3292 19848
rect 3424 19796 3476 19848
rect 3516 19796 3568 19848
rect 3976 19796 4028 19848
rect 12532 20000 12584 20052
rect 13452 20000 13504 20052
rect 15752 20043 15804 20052
rect 15752 20009 15761 20043
rect 15761 20009 15795 20043
rect 15795 20009 15804 20043
rect 15752 20000 15804 20009
rect 16212 20000 16264 20052
rect 16396 20043 16448 20052
rect 16396 20009 16405 20043
rect 16405 20009 16439 20043
rect 16439 20009 16448 20043
rect 16396 20000 16448 20009
rect 17408 20000 17460 20052
rect 20536 20000 20588 20052
rect 13360 19907 13412 19916
rect 13360 19873 13369 19907
rect 13369 19873 13403 19907
rect 13403 19873 13412 19907
rect 13360 19864 13412 19873
rect 20168 19932 20220 19984
rect 6736 19796 6788 19848
rect 12900 19796 12952 19848
rect 13084 19796 13136 19848
rect 13176 19839 13228 19848
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 13176 19796 13228 19805
rect 13268 19839 13320 19848
rect 13268 19805 13277 19839
rect 13277 19805 13311 19839
rect 13311 19805 13320 19839
rect 13268 19796 13320 19805
rect 15200 19796 15252 19848
rect 16304 19796 16356 19848
rect 17592 19839 17644 19848
rect 15384 19771 15436 19780
rect 15384 19737 15393 19771
rect 15393 19737 15427 19771
rect 15427 19737 15436 19771
rect 15384 19728 15436 19737
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 2964 19703 3016 19712
rect 2964 19669 2973 19703
rect 2973 19669 3007 19703
rect 3007 19669 3016 19703
rect 2964 19660 3016 19669
rect 3056 19660 3108 19712
rect 3424 19660 3476 19712
rect 4620 19660 4672 19712
rect 4804 19660 4856 19712
rect 16028 19660 16080 19712
rect 16764 19660 16816 19712
rect 18144 19660 18196 19712
rect 19248 19703 19300 19712
rect 19248 19669 19257 19703
rect 19257 19669 19291 19703
rect 19291 19669 19300 19703
rect 19248 19660 19300 19669
rect 20628 19660 20680 19712
rect 4255 19558 4307 19610
rect 4319 19558 4371 19610
rect 4383 19558 4435 19610
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 9545 19558 9597 19610
rect 9609 19558 9661 19610
rect 9673 19558 9725 19610
rect 9737 19558 9789 19610
rect 9801 19558 9853 19610
rect 14835 19558 14887 19610
rect 14899 19558 14951 19610
rect 14963 19558 15015 19610
rect 15027 19558 15079 19610
rect 15091 19558 15143 19610
rect 20125 19558 20177 19610
rect 20189 19558 20241 19610
rect 20253 19558 20305 19610
rect 20317 19558 20369 19610
rect 20381 19558 20433 19610
rect 2596 19388 2648 19440
rect 3332 19456 3384 19508
rect 3976 19456 4028 19508
rect 6828 19456 6880 19508
rect 8576 19456 8628 19508
rect 12900 19456 12952 19508
rect 3056 19363 3108 19372
rect 3056 19329 3065 19363
rect 3065 19329 3099 19363
rect 3099 19329 3108 19363
rect 3056 19320 3108 19329
rect 3240 19320 3292 19372
rect 3424 19320 3476 19372
rect 6000 19431 6052 19440
rect 6000 19397 6009 19431
rect 6009 19397 6043 19431
rect 6043 19397 6052 19431
rect 6000 19388 6052 19397
rect 5908 19363 5960 19372
rect 5908 19329 5917 19363
rect 5917 19329 5951 19363
rect 5951 19329 5960 19363
rect 5908 19320 5960 19329
rect 6184 19363 6236 19372
rect 6184 19329 6193 19363
rect 6193 19329 6227 19363
rect 6227 19329 6236 19363
rect 6184 19320 6236 19329
rect 6828 19363 6880 19372
rect 6828 19329 6837 19363
rect 6837 19329 6871 19363
rect 6871 19329 6880 19363
rect 6828 19320 6880 19329
rect 6276 19252 6328 19304
rect 9220 19320 9272 19372
rect 10416 19320 10468 19372
rect 12992 19388 13044 19440
rect 13268 19456 13320 19508
rect 16304 19456 16356 19508
rect 13360 19388 13412 19440
rect 17592 19456 17644 19508
rect 19248 19456 19300 19508
rect 8392 19295 8444 19304
rect 8392 19261 8401 19295
rect 8401 19261 8435 19295
rect 8435 19261 8444 19295
rect 8392 19252 8444 19261
rect 8668 19184 8720 19236
rect 11152 19320 11204 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 11980 19252 12032 19304
rect 13544 19320 13596 19372
rect 16304 19363 16356 19372
rect 16304 19329 16313 19363
rect 16313 19329 16347 19363
rect 16347 19329 16356 19363
rect 16304 19320 16356 19329
rect 16764 19363 16816 19372
rect 16764 19329 16773 19363
rect 16773 19329 16807 19363
rect 16807 19329 16816 19363
rect 16764 19320 16816 19329
rect 17408 19363 17460 19372
rect 16580 19252 16632 19304
rect 17408 19329 17417 19363
rect 17417 19329 17451 19363
rect 17451 19329 17460 19363
rect 17408 19320 17460 19329
rect 18328 19320 18380 19372
rect 19064 19363 19116 19372
rect 19064 19329 19073 19363
rect 19073 19329 19107 19363
rect 19107 19329 19116 19363
rect 19064 19320 19116 19329
rect 17040 19295 17092 19304
rect 17040 19261 17049 19295
rect 17049 19261 17083 19295
rect 17083 19261 17092 19295
rect 17040 19252 17092 19261
rect 19340 19252 19392 19304
rect 3332 19116 3384 19168
rect 3976 19116 4028 19168
rect 6552 19116 6604 19168
rect 6644 19116 6696 19168
rect 7196 19159 7248 19168
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 7472 19159 7524 19168
rect 7472 19125 7481 19159
rect 7481 19125 7515 19159
rect 7515 19125 7524 19159
rect 7472 19116 7524 19125
rect 7932 19159 7984 19168
rect 7932 19125 7941 19159
rect 7941 19125 7975 19159
rect 7975 19125 7984 19159
rect 7932 19116 7984 19125
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 10232 19116 10284 19168
rect 10876 19159 10928 19168
rect 10876 19125 10885 19159
rect 10885 19125 10919 19159
rect 10919 19125 10928 19159
rect 10876 19116 10928 19125
rect 12072 19116 12124 19168
rect 16212 19116 16264 19168
rect 17040 19116 17092 19168
rect 17132 19159 17184 19168
rect 17132 19125 17141 19159
rect 17141 19125 17175 19159
rect 17175 19125 17184 19159
rect 17132 19116 17184 19125
rect 19892 19116 19944 19168
rect 3595 19014 3647 19066
rect 3659 19014 3711 19066
rect 3723 19014 3775 19066
rect 3787 19014 3839 19066
rect 3851 19014 3903 19066
rect 8885 19014 8937 19066
rect 8949 19014 9001 19066
rect 9013 19014 9065 19066
rect 9077 19014 9129 19066
rect 9141 19014 9193 19066
rect 14175 19014 14227 19066
rect 14239 19014 14291 19066
rect 14303 19014 14355 19066
rect 14367 19014 14419 19066
rect 14431 19014 14483 19066
rect 19465 19014 19517 19066
rect 19529 19014 19581 19066
rect 19593 19014 19645 19066
rect 19657 19014 19709 19066
rect 19721 19014 19773 19066
rect 2596 18912 2648 18964
rect 4068 18912 4120 18964
rect 7656 18912 7708 18964
rect 9220 18955 9272 18964
rect 9220 18921 9229 18955
rect 9229 18921 9263 18955
rect 9263 18921 9272 18955
rect 9220 18912 9272 18921
rect 10876 18912 10928 18964
rect 11980 18912 12032 18964
rect 16304 18912 16356 18964
rect 16948 18912 17000 18964
rect 17132 18912 17184 18964
rect 17776 18912 17828 18964
rect 18328 18912 18380 18964
rect 4712 18819 4764 18828
rect 4712 18785 4721 18819
rect 4721 18785 4755 18819
rect 4755 18785 4764 18819
rect 4712 18776 4764 18785
rect 4896 18819 4948 18828
rect 4896 18785 4905 18819
rect 4905 18785 4939 18819
rect 4939 18785 4948 18819
rect 4896 18776 4948 18785
rect 6092 18776 6144 18828
rect 2780 18640 2832 18692
rect 3976 18572 4028 18624
rect 4160 18572 4212 18624
rect 4620 18708 4672 18760
rect 6736 18751 6788 18760
rect 6736 18717 6745 18751
rect 6745 18717 6779 18751
rect 6779 18717 6788 18751
rect 6736 18708 6788 18717
rect 6368 18640 6420 18692
rect 6644 18640 6696 18692
rect 4620 18572 4672 18624
rect 5540 18572 5592 18624
rect 6276 18615 6328 18624
rect 6276 18581 6285 18615
rect 6285 18581 6319 18615
rect 6319 18581 6328 18615
rect 6276 18572 6328 18581
rect 7196 18776 7248 18828
rect 8392 18776 8444 18828
rect 8852 18776 8904 18828
rect 7380 18751 7432 18760
rect 7380 18717 7389 18751
rect 7389 18717 7423 18751
rect 7423 18717 7432 18751
rect 7380 18708 7432 18717
rect 7932 18708 7984 18760
rect 9956 18708 10008 18760
rect 10232 18708 10284 18760
rect 11520 18708 11572 18760
rect 8300 18640 8352 18692
rect 8668 18640 8720 18692
rect 9220 18683 9272 18692
rect 9220 18649 9229 18683
rect 9229 18649 9263 18683
rect 9263 18649 9272 18683
rect 9220 18640 9272 18649
rect 11244 18640 11296 18692
rect 14096 18708 14148 18760
rect 16580 18844 16632 18896
rect 15568 18776 15620 18828
rect 18052 18776 18104 18828
rect 12440 18640 12492 18692
rect 12624 18640 12676 18692
rect 14372 18640 14424 18692
rect 14556 18640 14608 18692
rect 15200 18640 15252 18692
rect 8208 18572 8260 18624
rect 10232 18572 10284 18624
rect 11152 18572 11204 18624
rect 12072 18572 12124 18624
rect 12808 18572 12860 18624
rect 13544 18572 13596 18624
rect 17132 18640 17184 18692
rect 18144 18751 18196 18760
rect 18144 18717 18153 18751
rect 18153 18717 18187 18751
rect 18187 18717 18196 18751
rect 18144 18708 18196 18717
rect 19340 18708 19392 18760
rect 17500 18640 17552 18692
rect 19892 18640 19944 18692
rect 19248 18615 19300 18624
rect 19248 18581 19257 18615
rect 19257 18581 19291 18615
rect 19291 18581 19300 18615
rect 19248 18572 19300 18581
rect 4255 18470 4307 18522
rect 4319 18470 4371 18522
rect 4383 18470 4435 18522
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 9545 18470 9597 18522
rect 9609 18470 9661 18522
rect 9673 18470 9725 18522
rect 9737 18470 9789 18522
rect 9801 18470 9853 18522
rect 14835 18470 14887 18522
rect 14899 18470 14951 18522
rect 14963 18470 15015 18522
rect 15027 18470 15079 18522
rect 15091 18470 15143 18522
rect 20125 18470 20177 18522
rect 20189 18470 20241 18522
rect 20253 18470 20305 18522
rect 20317 18470 20369 18522
rect 20381 18470 20433 18522
rect 2780 18411 2832 18420
rect 2780 18377 2789 18411
rect 2789 18377 2823 18411
rect 2823 18377 2832 18411
rect 2780 18368 2832 18377
rect 4160 18411 4212 18420
rect 4160 18377 4169 18411
rect 4169 18377 4203 18411
rect 4203 18377 4212 18411
rect 4160 18368 4212 18377
rect 2964 18275 3016 18284
rect 2964 18241 2973 18275
rect 2973 18241 3007 18275
rect 3007 18241 3016 18275
rect 2964 18232 3016 18241
rect 4712 18368 4764 18420
rect 4804 18411 4856 18420
rect 4804 18377 4813 18411
rect 4813 18377 4847 18411
rect 4847 18377 4856 18411
rect 4804 18368 4856 18377
rect 5908 18368 5960 18420
rect 6368 18411 6420 18420
rect 6368 18377 6377 18411
rect 6377 18377 6411 18411
rect 6411 18377 6420 18411
rect 6368 18368 6420 18377
rect 7288 18368 7340 18420
rect 8852 18411 8904 18420
rect 8852 18377 8861 18411
rect 8861 18377 8895 18411
rect 8895 18377 8904 18411
rect 8852 18368 8904 18377
rect 11244 18411 11296 18420
rect 11244 18377 11253 18411
rect 11253 18377 11287 18411
rect 11287 18377 11296 18411
rect 11244 18368 11296 18377
rect 11520 18411 11572 18420
rect 11520 18377 11529 18411
rect 11529 18377 11563 18411
rect 11563 18377 11572 18411
rect 11520 18368 11572 18377
rect 11980 18368 12032 18420
rect 13176 18368 13228 18420
rect 14372 18411 14424 18420
rect 14372 18377 14381 18411
rect 14381 18377 14415 18411
rect 14415 18377 14424 18411
rect 14372 18368 14424 18377
rect 5080 18300 5132 18352
rect 11704 18300 11756 18352
rect 3976 18164 4028 18216
rect 4528 18275 4580 18284
rect 4528 18241 4537 18275
rect 4537 18241 4571 18275
rect 4571 18241 4580 18275
rect 4528 18232 4580 18241
rect 4712 18275 4764 18284
rect 4712 18241 4721 18275
rect 4721 18241 4755 18275
rect 4755 18241 4764 18275
rect 4712 18232 4764 18241
rect 3332 18028 3384 18080
rect 5540 18275 5592 18284
rect 5540 18241 5549 18275
rect 5549 18241 5583 18275
rect 5583 18241 5592 18275
rect 5540 18232 5592 18241
rect 5908 18232 5960 18284
rect 6092 18232 6144 18284
rect 6460 18232 6512 18284
rect 6552 18275 6604 18284
rect 6552 18241 6561 18275
rect 6561 18241 6595 18275
rect 6595 18241 6604 18275
rect 6552 18232 6604 18241
rect 6644 18232 6696 18284
rect 7472 18232 7524 18284
rect 5632 18207 5684 18216
rect 5632 18173 5641 18207
rect 5641 18173 5675 18207
rect 5675 18173 5684 18207
rect 5632 18164 5684 18173
rect 6000 18096 6052 18148
rect 6736 18028 6788 18080
rect 8208 18232 8260 18284
rect 10232 18232 10284 18284
rect 10876 18232 10928 18284
rect 11336 18275 11388 18284
rect 11336 18241 11345 18275
rect 11345 18241 11379 18275
rect 11379 18241 11388 18275
rect 11336 18232 11388 18241
rect 12624 18300 12676 18352
rect 12532 18275 12584 18284
rect 12532 18241 12541 18275
rect 12541 18241 12575 18275
rect 12575 18241 12584 18275
rect 12532 18232 12584 18241
rect 12992 18232 13044 18284
rect 13544 18232 13596 18284
rect 13728 18232 13780 18284
rect 8484 18164 8536 18216
rect 9680 18207 9732 18216
rect 9680 18173 9689 18207
rect 9689 18173 9723 18207
rect 9723 18173 9732 18207
rect 9680 18164 9732 18173
rect 8576 18096 8628 18148
rect 9220 18096 9272 18148
rect 12440 18164 12492 18216
rect 12808 18207 12860 18216
rect 12808 18173 12817 18207
rect 12817 18173 12851 18207
rect 12851 18173 12860 18207
rect 12808 18164 12860 18173
rect 14004 18207 14056 18216
rect 14004 18173 14013 18207
rect 14013 18173 14047 18207
rect 14047 18173 14056 18207
rect 14004 18164 14056 18173
rect 14740 18300 14792 18352
rect 14924 18300 14976 18352
rect 14648 18232 14700 18284
rect 14832 18207 14884 18216
rect 14832 18173 14841 18207
rect 14841 18173 14875 18207
rect 14875 18173 14884 18207
rect 15200 18343 15252 18352
rect 15200 18309 15209 18343
rect 15209 18309 15243 18343
rect 15243 18309 15252 18343
rect 17500 18343 17552 18352
rect 15200 18300 15252 18309
rect 17500 18309 17509 18343
rect 17509 18309 17543 18343
rect 17543 18309 17552 18343
rect 17500 18300 17552 18309
rect 14832 18164 14884 18173
rect 14648 18096 14700 18148
rect 17040 18164 17092 18216
rect 17132 18207 17184 18216
rect 17132 18173 17141 18207
rect 17141 18173 17175 18207
rect 17175 18173 17184 18207
rect 17132 18164 17184 18173
rect 8760 18028 8812 18080
rect 14556 18028 14608 18080
rect 14740 18071 14792 18080
rect 14740 18037 14749 18071
rect 14749 18037 14783 18071
rect 14783 18037 14792 18071
rect 14740 18028 14792 18037
rect 14924 18028 14976 18080
rect 16580 18028 16632 18080
rect 17040 18071 17092 18080
rect 17040 18037 17049 18071
rect 17049 18037 17083 18071
rect 17083 18037 17092 18071
rect 17040 18028 17092 18037
rect 3595 17926 3647 17978
rect 3659 17926 3711 17978
rect 3723 17926 3775 17978
rect 3787 17926 3839 17978
rect 3851 17926 3903 17978
rect 8885 17926 8937 17978
rect 8949 17926 9001 17978
rect 9013 17926 9065 17978
rect 9077 17926 9129 17978
rect 9141 17926 9193 17978
rect 14175 17926 14227 17978
rect 14239 17926 14291 17978
rect 14303 17926 14355 17978
rect 14367 17926 14419 17978
rect 14431 17926 14483 17978
rect 19465 17926 19517 17978
rect 19529 17926 19581 17978
rect 19593 17926 19645 17978
rect 19657 17926 19709 17978
rect 19721 17926 19773 17978
rect 9956 17824 10008 17876
rect 11336 17824 11388 17876
rect 12256 17824 12308 17876
rect 16028 17824 16080 17876
rect 17040 17824 17092 17876
rect 17408 17824 17460 17876
rect 4068 17688 4120 17740
rect 4528 17688 4580 17740
rect 3332 17620 3384 17672
rect 3516 17620 3568 17672
rect 5540 17620 5592 17672
rect 9312 17620 9364 17672
rect 10048 17663 10100 17672
rect 10048 17629 10057 17663
rect 10057 17629 10091 17663
rect 10091 17629 10100 17663
rect 10048 17620 10100 17629
rect 13728 17756 13780 17808
rect 10324 17595 10376 17604
rect 10324 17561 10333 17595
rect 10333 17561 10367 17595
rect 10367 17561 10376 17595
rect 10324 17552 10376 17561
rect 11336 17620 11388 17672
rect 11888 17663 11940 17672
rect 11888 17629 11897 17663
rect 11897 17629 11931 17663
rect 11931 17629 11940 17663
rect 11888 17620 11940 17629
rect 12072 17620 12124 17672
rect 12624 17663 12676 17672
rect 12624 17629 12633 17663
rect 12633 17629 12667 17663
rect 12667 17629 12676 17663
rect 12624 17620 12676 17629
rect 13452 17620 13504 17672
rect 14832 17688 14884 17740
rect 15292 17620 15344 17672
rect 3516 17527 3568 17536
rect 3516 17493 3525 17527
rect 3525 17493 3559 17527
rect 3559 17493 3568 17527
rect 3516 17484 3568 17493
rect 3792 17527 3844 17536
rect 3792 17493 3801 17527
rect 3801 17493 3835 17527
rect 3835 17493 3844 17527
rect 3792 17484 3844 17493
rect 4160 17484 4212 17536
rect 4712 17484 4764 17536
rect 5172 17484 5224 17536
rect 9312 17484 9364 17536
rect 10140 17527 10192 17536
rect 10140 17493 10149 17527
rect 10149 17493 10183 17527
rect 10183 17493 10192 17527
rect 10140 17484 10192 17493
rect 12440 17527 12492 17536
rect 12440 17493 12449 17527
rect 12449 17493 12483 17527
rect 12483 17493 12492 17527
rect 12440 17484 12492 17493
rect 13268 17552 13320 17604
rect 14556 17552 14608 17604
rect 16212 17663 16264 17672
rect 16212 17629 16221 17663
rect 16221 17629 16255 17663
rect 16255 17629 16264 17663
rect 16212 17620 16264 17629
rect 16580 17663 16632 17672
rect 16580 17629 16614 17663
rect 16614 17629 16632 17663
rect 16580 17620 16632 17629
rect 16948 17620 17000 17672
rect 19800 17620 19852 17672
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 12992 17484 13044 17536
rect 14648 17484 14700 17536
rect 15568 17484 15620 17536
rect 19892 17527 19944 17536
rect 19892 17493 19901 17527
rect 19901 17493 19935 17527
rect 19935 17493 19944 17527
rect 19892 17484 19944 17493
rect 20904 17527 20956 17536
rect 20904 17493 20913 17527
rect 20913 17493 20947 17527
rect 20947 17493 20956 17527
rect 20904 17484 20956 17493
rect 4255 17382 4307 17434
rect 4319 17382 4371 17434
rect 4383 17382 4435 17434
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 9545 17382 9597 17434
rect 9609 17382 9661 17434
rect 9673 17382 9725 17434
rect 9737 17382 9789 17434
rect 9801 17382 9853 17434
rect 14835 17382 14887 17434
rect 14899 17382 14951 17434
rect 14963 17382 15015 17434
rect 15027 17382 15079 17434
rect 15091 17382 15143 17434
rect 20125 17382 20177 17434
rect 20189 17382 20241 17434
rect 20253 17382 20305 17434
rect 20317 17382 20369 17434
rect 20381 17382 20433 17434
rect 3516 17280 3568 17332
rect 3792 17280 3844 17332
rect 4620 17280 4672 17332
rect 10324 17280 10376 17332
rect 12532 17280 12584 17332
rect 14648 17280 14700 17332
rect 14740 17280 14792 17332
rect 19892 17280 19944 17332
rect 21456 17280 21508 17332
rect 1492 17144 1544 17196
rect 3608 17187 3660 17196
rect 3608 17153 3617 17187
rect 3617 17153 3651 17187
rect 3651 17153 3660 17187
rect 3608 17144 3660 17153
rect 6184 17212 6236 17264
rect 9496 17212 9548 17264
rect 13912 17212 13964 17264
rect 14556 17212 14608 17264
rect 4160 17144 4212 17196
rect 4436 17187 4488 17196
rect 4436 17153 4445 17187
rect 4445 17153 4479 17187
rect 4479 17153 4488 17187
rect 4436 17144 4488 17153
rect 4712 17144 4764 17196
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 6644 17187 6696 17196
rect 6644 17153 6653 17187
rect 6653 17153 6687 17187
rect 6687 17153 6696 17187
rect 6644 17144 6696 17153
rect 7288 17187 7340 17196
rect 7288 17153 7297 17187
rect 7297 17153 7331 17187
rect 7331 17153 7340 17187
rect 7288 17144 7340 17153
rect 7840 17144 7892 17196
rect 9312 17187 9364 17196
rect 9312 17153 9335 17187
rect 9335 17153 9364 17187
rect 4068 17008 4120 17060
rect 7104 17076 7156 17128
rect 8208 17008 8260 17060
rect 9312 17144 9364 17153
rect 8576 17076 8628 17128
rect 3240 16983 3292 16992
rect 3240 16949 3249 16983
rect 3249 16949 3283 16983
rect 3283 16949 3292 16983
rect 3240 16940 3292 16949
rect 5264 16940 5316 16992
rect 6092 16940 6144 16992
rect 7472 16983 7524 16992
rect 7472 16949 7481 16983
rect 7481 16949 7515 16983
rect 7515 16949 7524 16983
rect 7472 16940 7524 16949
rect 7564 16983 7616 16992
rect 7564 16949 7573 16983
rect 7573 16949 7607 16983
rect 7607 16949 7616 16983
rect 7564 16940 7616 16949
rect 8484 16940 8536 16992
rect 11244 17119 11296 17128
rect 11244 17085 11253 17119
rect 11253 17085 11287 17119
rect 11287 17085 11296 17119
rect 11244 17076 11296 17085
rect 12256 17076 12308 17128
rect 12532 17076 12584 17128
rect 12808 17187 12860 17196
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 12900 17187 12952 17196
rect 12900 17153 12909 17187
rect 12909 17153 12943 17187
rect 12943 17153 12952 17187
rect 12900 17144 12952 17153
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 15568 17255 15620 17264
rect 15568 17221 15577 17255
rect 15577 17221 15611 17255
rect 15611 17221 15620 17255
rect 15568 17212 15620 17221
rect 15292 17144 15344 17196
rect 15476 17144 15528 17196
rect 16212 17144 16264 17196
rect 9404 16940 9456 16992
rect 10048 16940 10100 16992
rect 11336 16940 11388 16992
rect 11612 16940 11664 16992
rect 15200 17008 15252 17060
rect 16948 17076 17000 17128
rect 19340 17212 19392 17264
rect 18512 17144 18564 17196
rect 19892 17187 19944 17196
rect 19892 17153 19901 17187
rect 19901 17153 19935 17187
rect 19935 17153 19944 17187
rect 19892 17144 19944 17153
rect 12992 16940 13044 16992
rect 13360 16983 13412 16992
rect 13360 16949 13369 16983
rect 13369 16949 13403 16983
rect 13403 16949 13412 16983
rect 13360 16940 13412 16949
rect 20076 16940 20128 16992
rect 3595 16838 3647 16890
rect 3659 16838 3711 16890
rect 3723 16838 3775 16890
rect 3787 16838 3839 16890
rect 3851 16838 3903 16890
rect 8885 16838 8937 16890
rect 8949 16838 9001 16890
rect 9013 16838 9065 16890
rect 9077 16838 9129 16890
rect 9141 16838 9193 16890
rect 14175 16838 14227 16890
rect 14239 16838 14291 16890
rect 14303 16838 14355 16890
rect 14367 16838 14419 16890
rect 14431 16838 14483 16890
rect 19465 16838 19517 16890
rect 19529 16838 19581 16890
rect 19593 16838 19645 16890
rect 19657 16838 19709 16890
rect 19721 16838 19773 16890
rect 3332 16668 3384 16720
rect 1492 16600 1544 16652
rect 4896 16736 4948 16788
rect 5632 16736 5684 16788
rect 6368 16736 6420 16788
rect 6460 16779 6512 16788
rect 6460 16745 6469 16779
rect 6469 16745 6503 16779
rect 6503 16745 6512 16779
rect 6460 16736 6512 16745
rect 7104 16668 7156 16720
rect 4620 16643 4672 16652
rect 4620 16609 4629 16643
rect 4629 16609 4663 16643
rect 4663 16609 4672 16643
rect 4620 16600 4672 16609
rect 6552 16600 6604 16652
rect 3516 16532 3568 16584
rect 4436 16575 4488 16584
rect 4436 16541 4445 16575
rect 4445 16541 4479 16575
rect 4479 16541 4488 16575
rect 4436 16532 4488 16541
rect 2136 16464 2188 16516
rect 4068 16464 4120 16516
rect 6920 16575 6972 16584
rect 6920 16541 6929 16575
rect 6929 16541 6963 16575
rect 6963 16541 6972 16575
rect 6920 16532 6972 16541
rect 7380 16736 7432 16788
rect 8208 16668 8260 16720
rect 7472 16575 7524 16584
rect 7472 16541 7506 16575
rect 7506 16541 7524 16575
rect 7472 16532 7524 16541
rect 5724 16464 5776 16516
rect 12072 16736 12124 16788
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 12900 16779 12952 16788
rect 12900 16745 12909 16779
rect 12909 16745 12943 16779
rect 12943 16745 12952 16779
rect 12900 16736 12952 16745
rect 14648 16736 14700 16788
rect 15292 16736 15344 16788
rect 18512 16736 18564 16788
rect 19800 16736 19852 16788
rect 20904 16736 20956 16788
rect 11244 16711 11296 16720
rect 11244 16677 11253 16711
rect 11253 16677 11287 16711
rect 11287 16677 11296 16711
rect 11244 16668 11296 16677
rect 12624 16668 12676 16720
rect 9404 16600 9456 16652
rect 9496 16575 9548 16584
rect 9496 16541 9505 16575
rect 9505 16541 9539 16575
rect 9539 16541 9548 16575
rect 9496 16532 9548 16541
rect 9772 16575 9824 16584
rect 9772 16541 9781 16575
rect 9781 16541 9815 16575
rect 9815 16541 9824 16575
rect 9772 16532 9824 16541
rect 12440 16600 12492 16652
rect 11336 16532 11388 16584
rect 13268 16600 13320 16652
rect 15476 16600 15528 16652
rect 18328 16600 18380 16652
rect 19248 16600 19300 16652
rect 20076 16600 20128 16652
rect 1676 16396 1728 16448
rect 3516 16396 3568 16448
rect 4804 16396 4856 16448
rect 8484 16464 8536 16516
rect 7472 16396 7524 16448
rect 8576 16439 8628 16448
rect 8576 16405 8585 16439
rect 8585 16405 8619 16439
rect 8619 16405 8628 16439
rect 12716 16532 12768 16584
rect 8576 16396 8628 16405
rect 11428 16396 11480 16448
rect 12348 16396 12400 16448
rect 12992 16464 13044 16516
rect 13176 16575 13228 16584
rect 13176 16541 13185 16575
rect 13185 16541 13219 16575
rect 13219 16541 13228 16575
rect 13176 16532 13228 16541
rect 13452 16575 13504 16584
rect 13452 16541 13461 16575
rect 13461 16541 13495 16575
rect 13495 16541 13504 16575
rect 13452 16532 13504 16541
rect 15568 16575 15620 16584
rect 15568 16541 15577 16575
rect 15577 16541 15611 16575
rect 15611 16541 15620 16575
rect 15568 16532 15620 16541
rect 17592 16575 17644 16584
rect 17592 16541 17601 16575
rect 17601 16541 17635 16575
rect 17635 16541 17644 16575
rect 17592 16532 17644 16541
rect 13360 16464 13412 16516
rect 19064 16575 19116 16584
rect 19064 16541 19073 16575
rect 19073 16541 19107 16575
rect 19107 16541 19116 16575
rect 19064 16532 19116 16541
rect 21640 16575 21692 16584
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 12808 16396 12860 16448
rect 14464 16396 14516 16448
rect 14740 16396 14792 16448
rect 17224 16396 17276 16448
rect 18052 16396 18104 16448
rect 19708 16396 19760 16448
rect 19984 16396 20036 16448
rect 20720 16396 20772 16448
rect 4255 16294 4307 16346
rect 4319 16294 4371 16346
rect 4383 16294 4435 16346
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 9545 16294 9597 16346
rect 9609 16294 9661 16346
rect 9673 16294 9725 16346
rect 9737 16294 9789 16346
rect 9801 16294 9853 16346
rect 14835 16294 14887 16346
rect 14899 16294 14951 16346
rect 14963 16294 15015 16346
rect 15027 16294 15079 16346
rect 15091 16294 15143 16346
rect 20125 16294 20177 16346
rect 20189 16294 20241 16346
rect 20253 16294 20305 16346
rect 20317 16294 20369 16346
rect 20381 16294 20433 16346
rect 1676 16192 1728 16244
rect 4620 16192 4672 16244
rect 5724 16235 5776 16244
rect 5724 16201 5733 16235
rect 5733 16201 5767 16235
rect 5767 16201 5776 16235
rect 5724 16192 5776 16201
rect 6920 16192 6972 16244
rect 8300 16235 8352 16244
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 8300 16192 8352 16201
rect 9404 16192 9456 16244
rect 2136 16124 2188 16176
rect 11796 16192 11848 16244
rect 11428 16124 11480 16176
rect 11612 16167 11664 16176
rect 11612 16133 11621 16167
rect 11621 16133 11655 16167
rect 11655 16133 11664 16167
rect 11612 16124 11664 16133
rect 2320 16099 2372 16108
rect 2320 16065 2329 16099
rect 2329 16065 2363 16099
rect 2363 16065 2372 16099
rect 2320 16056 2372 16065
rect 3240 16056 3292 16108
rect 4528 16056 4580 16108
rect 4804 16099 4856 16108
rect 4804 16065 4813 16099
rect 4813 16065 4847 16099
rect 4847 16065 4856 16099
rect 4804 16056 4856 16065
rect 5264 16099 5316 16108
rect 5264 16065 5273 16099
rect 5273 16065 5307 16099
rect 5307 16065 5316 16099
rect 5264 16056 5316 16065
rect 5356 16056 5408 16108
rect 6092 16056 6144 16108
rect 6368 16099 6420 16108
rect 6368 16065 6377 16099
rect 6377 16065 6411 16099
rect 6411 16065 6420 16099
rect 6368 16056 6420 16065
rect 6460 16056 6512 16108
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 7104 16056 7156 16108
rect 7472 16099 7524 16108
rect 7472 16065 7481 16099
rect 7481 16065 7515 16099
rect 7515 16065 7524 16099
rect 7472 16056 7524 16065
rect 5540 15988 5592 16040
rect 4620 15852 4672 15904
rect 4988 15895 5040 15904
rect 4988 15861 4997 15895
rect 4997 15861 5031 15895
rect 5031 15861 5040 15895
rect 4988 15852 5040 15861
rect 7656 16056 7708 16108
rect 8208 16056 8260 16108
rect 9220 16056 9272 16108
rect 10324 16056 10376 16108
rect 11336 16031 11388 16040
rect 11336 15997 11345 16031
rect 11345 15997 11379 16031
rect 11379 15997 11388 16031
rect 11336 15988 11388 15997
rect 11520 16099 11572 16108
rect 11520 16065 11529 16099
rect 11529 16065 11563 16099
rect 11563 16065 11572 16099
rect 11520 16056 11572 16065
rect 15200 16192 15252 16244
rect 15476 16192 15528 16244
rect 19064 16235 19116 16244
rect 19064 16201 19073 16235
rect 19073 16201 19107 16235
rect 19107 16201 19116 16235
rect 19064 16192 19116 16201
rect 19800 16192 19852 16244
rect 19984 16192 20036 16244
rect 12624 16124 12676 16176
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 12808 16099 12860 16108
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 14556 16124 14608 16176
rect 6644 15920 6696 15972
rect 13268 15988 13320 16040
rect 11888 15920 11940 15972
rect 12072 15963 12124 15972
rect 12072 15929 12081 15963
rect 12081 15929 12115 15963
rect 12115 15929 12124 15963
rect 12072 15920 12124 15929
rect 12440 15920 12492 15972
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 14648 16056 14700 16108
rect 14096 15988 14148 16040
rect 14924 16056 14976 16108
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 17224 16099 17276 16108
rect 17224 16065 17258 16099
rect 17258 16065 17276 16099
rect 17224 16056 17276 16065
rect 19616 15920 19668 15972
rect 19892 16056 19944 16108
rect 20352 16192 20404 16244
rect 21456 16192 21508 16244
rect 21640 16235 21692 16244
rect 21640 16201 21649 16235
rect 21649 16201 21683 16235
rect 21683 16201 21692 16235
rect 21640 16192 21692 16201
rect 6552 15852 6604 15904
rect 10140 15852 10192 15904
rect 12256 15895 12308 15904
rect 12256 15861 12265 15895
rect 12265 15861 12299 15895
rect 12299 15861 12308 15895
rect 12256 15852 12308 15861
rect 14832 15852 14884 15904
rect 18420 15852 18472 15904
rect 19432 15852 19484 15904
rect 19708 15852 19760 15904
rect 19892 15852 19944 15904
rect 20260 15852 20312 15904
rect 3595 15750 3647 15802
rect 3659 15750 3711 15802
rect 3723 15750 3775 15802
rect 3787 15750 3839 15802
rect 3851 15750 3903 15802
rect 8885 15750 8937 15802
rect 8949 15750 9001 15802
rect 9013 15750 9065 15802
rect 9077 15750 9129 15802
rect 9141 15750 9193 15802
rect 14175 15750 14227 15802
rect 14239 15750 14291 15802
rect 14303 15750 14355 15802
rect 14367 15750 14419 15802
rect 14431 15750 14483 15802
rect 19465 15750 19517 15802
rect 19529 15750 19581 15802
rect 19593 15750 19645 15802
rect 19657 15750 19709 15802
rect 19721 15750 19773 15802
rect 2320 15691 2372 15700
rect 2320 15657 2329 15691
rect 2329 15657 2363 15691
rect 2363 15657 2372 15691
rect 2320 15648 2372 15657
rect 3240 15648 3292 15700
rect 3516 15648 3568 15700
rect 4712 15648 4764 15700
rect 4988 15648 5040 15700
rect 7288 15648 7340 15700
rect 7840 15691 7892 15700
rect 7840 15657 7849 15691
rect 7849 15657 7883 15691
rect 7883 15657 7892 15691
rect 7840 15648 7892 15657
rect 11796 15648 11848 15700
rect 12900 15648 12952 15700
rect 14556 15648 14608 15700
rect 16948 15691 17000 15700
rect 16948 15657 16957 15691
rect 16957 15657 16991 15691
rect 16991 15657 17000 15691
rect 16948 15648 17000 15657
rect 4068 15512 4120 15564
rect 4528 15512 4580 15564
rect 4620 15444 4672 15496
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 8576 15580 8628 15632
rect 8392 15512 8444 15564
rect 9220 15512 9272 15564
rect 12348 15512 12400 15564
rect 13820 15580 13872 15632
rect 19432 15648 19484 15700
rect 19984 15648 20036 15700
rect 20260 15691 20312 15700
rect 20260 15657 20269 15691
rect 20269 15657 20303 15691
rect 20303 15657 20312 15691
rect 20260 15648 20312 15657
rect 7564 15444 7616 15496
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 2596 15351 2648 15360
rect 2596 15317 2605 15351
rect 2605 15317 2639 15351
rect 2639 15317 2648 15351
rect 2596 15308 2648 15317
rect 3424 15376 3476 15428
rect 3056 15308 3108 15360
rect 4160 15308 4212 15360
rect 4712 15308 4764 15360
rect 4896 15351 4948 15360
rect 4896 15317 4905 15351
rect 4905 15317 4939 15351
rect 4939 15317 4948 15351
rect 4896 15308 4948 15317
rect 7472 15308 7524 15360
rect 7656 15308 7708 15360
rect 12164 15444 12216 15496
rect 12992 15512 13044 15564
rect 14280 15444 14332 15496
rect 14832 15444 14884 15496
rect 12808 15351 12860 15360
rect 12808 15317 12817 15351
rect 12817 15317 12851 15351
rect 12851 15317 12860 15351
rect 12808 15308 12860 15317
rect 13084 15308 13136 15360
rect 14924 15376 14976 15428
rect 15200 15487 15252 15496
rect 15200 15453 15209 15487
rect 15209 15453 15243 15487
rect 15243 15453 15252 15487
rect 15200 15444 15252 15453
rect 15292 15487 15344 15496
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 16672 15444 16724 15496
rect 18236 15487 18288 15496
rect 18236 15453 18245 15487
rect 18245 15453 18279 15487
rect 18279 15453 18288 15487
rect 18236 15444 18288 15453
rect 18420 15487 18472 15496
rect 18420 15453 18429 15487
rect 18429 15453 18463 15487
rect 18463 15453 18472 15487
rect 18420 15444 18472 15453
rect 19064 15487 19116 15496
rect 19064 15453 19073 15487
rect 19073 15453 19107 15487
rect 19107 15453 19116 15487
rect 19064 15444 19116 15453
rect 19892 15580 19944 15632
rect 15752 15376 15804 15428
rect 17592 15376 17644 15428
rect 19892 15444 19944 15496
rect 19616 15376 19668 15428
rect 19708 15376 19760 15428
rect 20352 15376 20404 15428
rect 20536 15487 20588 15496
rect 20536 15453 20545 15487
rect 20545 15453 20579 15487
rect 20579 15453 20588 15487
rect 20536 15444 20588 15453
rect 21640 15444 21692 15496
rect 20904 15376 20956 15428
rect 18328 15308 18380 15360
rect 18604 15351 18656 15360
rect 18604 15317 18613 15351
rect 18613 15317 18647 15351
rect 18647 15317 18656 15351
rect 18604 15308 18656 15317
rect 18880 15351 18932 15360
rect 18880 15317 18889 15351
rect 18889 15317 18923 15351
rect 18923 15317 18932 15351
rect 18880 15308 18932 15317
rect 19432 15308 19484 15360
rect 4255 15206 4307 15258
rect 4319 15206 4371 15258
rect 4383 15206 4435 15258
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 9545 15206 9597 15258
rect 9609 15206 9661 15258
rect 9673 15206 9725 15258
rect 9737 15206 9789 15258
rect 9801 15206 9853 15258
rect 14835 15206 14887 15258
rect 14899 15206 14951 15258
rect 14963 15206 15015 15258
rect 15027 15206 15079 15258
rect 15091 15206 15143 15258
rect 20125 15206 20177 15258
rect 20189 15206 20241 15258
rect 20253 15206 20305 15258
rect 20317 15206 20369 15258
rect 20381 15206 20433 15258
rect 2596 15036 2648 15088
rect 4160 15104 4212 15156
rect 4988 15104 5040 15156
rect 3516 15036 3568 15088
rect 4068 15036 4120 15088
rect 6552 15036 6604 15088
rect 8484 15036 8536 15088
rect 1492 14968 1544 15020
rect 3148 14900 3200 14952
rect 3424 14832 3476 14884
rect 4068 14943 4120 14952
rect 4068 14909 4077 14943
rect 4077 14909 4111 14943
rect 4111 14909 4120 14943
rect 4068 14900 4120 14909
rect 4252 14943 4304 14952
rect 4252 14909 4261 14943
rect 4261 14909 4295 14943
rect 4295 14909 4304 14943
rect 4252 14900 4304 14909
rect 4436 15011 4488 15020
rect 4436 14977 4445 15011
rect 4445 14977 4479 15011
rect 4479 14977 4488 15011
rect 4436 14968 4488 14977
rect 4528 15011 4580 15020
rect 4528 14977 4537 15011
rect 4537 14977 4571 15011
rect 4571 14977 4580 15011
rect 4528 14968 4580 14977
rect 4620 14900 4672 14952
rect 3332 14807 3384 14816
rect 3332 14773 3341 14807
rect 3341 14773 3375 14807
rect 3375 14773 3384 14807
rect 3332 14764 3384 14773
rect 3976 14807 4028 14816
rect 3976 14773 3985 14807
rect 3985 14773 4019 14807
rect 4019 14773 4028 14807
rect 3976 14764 4028 14773
rect 4712 14832 4764 14884
rect 6736 14968 6788 15020
rect 8392 14968 8444 15020
rect 12808 15104 12860 15156
rect 13820 15147 13872 15156
rect 13820 15113 13829 15147
rect 13829 15113 13863 15147
rect 13863 15113 13872 15147
rect 13820 15104 13872 15113
rect 14280 15104 14332 15156
rect 14648 15104 14700 15156
rect 15568 15104 15620 15156
rect 16672 15147 16724 15156
rect 16672 15113 16681 15147
rect 16681 15113 16715 15147
rect 16715 15113 16724 15147
rect 16672 15104 16724 15113
rect 14096 15036 14148 15088
rect 15200 14968 15252 15020
rect 15568 15011 15620 15020
rect 15568 14977 15577 15011
rect 15577 14977 15611 15011
rect 15611 14977 15620 15011
rect 15568 14968 15620 14977
rect 16948 14968 17000 15020
rect 18880 15104 18932 15156
rect 19708 15104 19760 15156
rect 19800 15147 19852 15156
rect 19800 15113 19809 15147
rect 19809 15113 19843 15147
rect 19843 15113 19852 15147
rect 19800 15104 19852 15113
rect 18604 15036 18656 15088
rect 18328 14968 18380 15020
rect 19340 15036 19392 15088
rect 7012 14832 7064 14884
rect 7656 14832 7708 14884
rect 18236 14900 18288 14952
rect 19432 14968 19484 15020
rect 19248 14832 19300 14884
rect 19892 14900 19944 14952
rect 20720 15104 20772 15156
rect 20904 15147 20956 15156
rect 20904 15113 20913 15147
rect 20913 15113 20947 15147
rect 20947 15113 20956 15147
rect 20904 15104 20956 15113
rect 19616 14832 19668 14884
rect 4160 14764 4212 14816
rect 5080 14764 5132 14816
rect 5816 14764 5868 14816
rect 6828 14764 6880 14816
rect 7380 14764 7432 14816
rect 14556 14764 14608 14816
rect 18420 14807 18472 14816
rect 18420 14773 18429 14807
rect 18429 14773 18463 14807
rect 18463 14773 18472 14807
rect 18420 14764 18472 14773
rect 19340 14764 19392 14816
rect 19892 14764 19944 14816
rect 19984 14807 20036 14816
rect 19984 14773 19993 14807
rect 19993 14773 20027 14807
rect 20027 14773 20036 14807
rect 19984 14764 20036 14773
rect 3595 14662 3647 14714
rect 3659 14662 3711 14714
rect 3723 14662 3775 14714
rect 3787 14662 3839 14714
rect 3851 14662 3903 14714
rect 8885 14662 8937 14714
rect 8949 14662 9001 14714
rect 9013 14662 9065 14714
rect 9077 14662 9129 14714
rect 9141 14662 9193 14714
rect 14175 14662 14227 14714
rect 14239 14662 14291 14714
rect 14303 14662 14355 14714
rect 14367 14662 14419 14714
rect 14431 14662 14483 14714
rect 19465 14662 19517 14714
rect 19529 14662 19581 14714
rect 19593 14662 19645 14714
rect 19657 14662 19709 14714
rect 19721 14662 19773 14714
rect 3148 14560 3200 14612
rect 3332 14560 3384 14612
rect 1492 14424 1544 14476
rect 4068 14560 4120 14612
rect 4436 14560 4488 14612
rect 4896 14560 4948 14612
rect 7472 14560 7524 14612
rect 8484 14560 8536 14612
rect 4528 14424 4580 14476
rect 5448 14424 5500 14476
rect 6000 14535 6052 14544
rect 6000 14501 6009 14535
rect 6009 14501 6043 14535
rect 6043 14501 6052 14535
rect 6000 14492 6052 14501
rect 8668 14535 8720 14544
rect 8668 14501 8677 14535
rect 8677 14501 8711 14535
rect 8711 14501 8720 14535
rect 8668 14492 8720 14501
rect 8760 14492 8812 14544
rect 3516 14356 3568 14408
rect 5080 14356 5132 14408
rect 3976 14288 4028 14340
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 6736 14356 6788 14365
rect 7012 14399 7064 14408
rect 7012 14365 7021 14399
rect 7021 14365 7055 14399
rect 7055 14365 7064 14399
rect 7012 14356 7064 14365
rect 6920 14331 6972 14340
rect 6920 14297 6929 14331
rect 6929 14297 6963 14331
rect 6963 14297 6972 14331
rect 7472 14399 7524 14408
rect 7472 14365 7481 14399
rect 7481 14365 7515 14399
rect 7515 14365 7524 14399
rect 7472 14356 7524 14365
rect 7840 14424 7892 14476
rect 9220 14492 9272 14544
rect 8024 14399 8076 14408
rect 8024 14365 8033 14399
rect 8033 14365 8067 14399
rect 8067 14365 8076 14399
rect 8024 14356 8076 14365
rect 8392 14356 8444 14408
rect 6920 14288 6972 14297
rect 9496 14399 9548 14408
rect 9496 14365 9505 14399
rect 9505 14365 9539 14399
rect 9539 14365 9548 14399
rect 9496 14356 9548 14365
rect 9312 14288 9364 14340
rect 10140 14356 10192 14408
rect 10232 14356 10284 14408
rect 10968 14356 11020 14408
rect 11888 14356 11940 14408
rect 12164 14356 12216 14408
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 14556 14603 14608 14612
rect 14556 14569 14565 14603
rect 14565 14569 14599 14603
rect 14599 14569 14608 14603
rect 14556 14560 14608 14569
rect 13728 14424 13780 14476
rect 15200 14603 15252 14612
rect 15200 14569 15209 14603
rect 15209 14569 15243 14603
rect 15243 14569 15252 14603
rect 15200 14560 15252 14569
rect 13084 14356 13136 14365
rect 15292 14424 15344 14476
rect 14648 14356 14700 14408
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 16304 14492 16356 14544
rect 18052 14560 18104 14612
rect 18604 14560 18656 14612
rect 16948 14424 17000 14476
rect 16764 14399 16816 14408
rect 16764 14365 16773 14399
rect 16773 14365 16807 14399
rect 16807 14365 16816 14399
rect 16764 14356 16816 14365
rect 19248 14560 19300 14612
rect 19340 14560 19392 14612
rect 7748 14220 7800 14272
rect 8392 14220 8444 14272
rect 8484 14220 8536 14272
rect 10048 14220 10100 14272
rect 10876 14263 10928 14272
rect 10876 14229 10885 14263
rect 10885 14229 10919 14263
rect 10919 14229 10928 14263
rect 10876 14220 10928 14229
rect 11612 14220 11664 14272
rect 12624 14263 12676 14272
rect 12624 14229 12633 14263
rect 12633 14229 12667 14263
rect 12667 14229 12676 14263
rect 12624 14220 12676 14229
rect 14372 14220 14424 14272
rect 14464 14220 14516 14272
rect 16948 14263 17000 14272
rect 16948 14229 16957 14263
rect 16957 14229 16991 14263
rect 16991 14229 17000 14263
rect 16948 14220 17000 14229
rect 17592 14288 17644 14340
rect 4255 14118 4307 14170
rect 4319 14118 4371 14170
rect 4383 14118 4435 14170
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 9545 14118 9597 14170
rect 9609 14118 9661 14170
rect 9673 14118 9725 14170
rect 9737 14118 9789 14170
rect 9801 14118 9853 14170
rect 14835 14118 14887 14170
rect 14899 14118 14951 14170
rect 14963 14118 15015 14170
rect 15027 14118 15079 14170
rect 15091 14118 15143 14170
rect 20125 14118 20177 14170
rect 20189 14118 20241 14170
rect 20253 14118 20305 14170
rect 20317 14118 20369 14170
rect 20381 14118 20433 14170
rect 3148 13923 3200 13932
rect 3148 13889 3157 13923
rect 3157 13889 3191 13923
rect 3191 13889 3200 13923
rect 3148 13880 3200 13889
rect 3976 14016 4028 14068
rect 4160 14016 4212 14068
rect 5448 14016 5500 14068
rect 5632 14016 5684 14068
rect 6736 14016 6788 14068
rect 8024 14016 8076 14068
rect 4344 13948 4396 14000
rect 5080 13948 5132 14000
rect 5172 13923 5224 13932
rect 5172 13889 5181 13923
rect 5181 13889 5215 13923
rect 5215 13889 5224 13923
rect 5172 13880 5224 13889
rect 5540 13880 5592 13932
rect 8484 14059 8536 14068
rect 8484 14025 8493 14059
rect 8493 14025 8527 14059
rect 8527 14025 8536 14059
rect 8484 14016 8536 14025
rect 8668 14016 8720 14068
rect 6644 13923 6696 13932
rect 6644 13889 6653 13923
rect 6653 13889 6687 13923
rect 6687 13889 6696 13923
rect 6644 13880 6696 13889
rect 7012 13880 7064 13932
rect 7380 13923 7432 13932
rect 7380 13889 7414 13923
rect 7414 13889 7432 13923
rect 7380 13880 7432 13889
rect 8300 13880 8352 13932
rect 8392 13880 8444 13932
rect 10232 14016 10284 14068
rect 10876 14016 10928 14068
rect 10968 14016 11020 14068
rect 5816 13855 5868 13864
rect 5816 13821 5825 13855
rect 5825 13821 5859 13855
rect 5859 13821 5868 13855
rect 5816 13812 5868 13821
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 10048 13880 10100 13932
rect 10784 13880 10836 13932
rect 12624 14016 12676 14068
rect 13176 14016 13228 14068
rect 13728 14016 13780 14068
rect 14372 14059 14424 14068
rect 14372 14025 14381 14059
rect 14381 14025 14415 14059
rect 14415 14025 14424 14059
rect 14372 14016 14424 14025
rect 14464 14016 14516 14068
rect 15200 14016 15252 14068
rect 15292 14016 15344 14068
rect 15384 14059 15436 14068
rect 15384 14025 15393 14059
rect 15393 14025 15427 14059
rect 15427 14025 15436 14059
rect 15384 14016 15436 14025
rect 15568 14016 15620 14068
rect 16304 14016 16356 14068
rect 16948 14016 17000 14068
rect 19064 14016 19116 14068
rect 15292 13880 15344 13932
rect 11336 13855 11388 13864
rect 11336 13821 11345 13855
rect 11345 13821 11379 13855
rect 11379 13821 11388 13855
rect 11336 13812 11388 13821
rect 11612 13812 11664 13864
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 15568 13812 15620 13864
rect 16764 13880 16816 13932
rect 18604 13880 18656 13932
rect 19984 13923 20036 13932
rect 19984 13889 19993 13923
rect 19993 13889 20027 13923
rect 20027 13889 20036 13923
rect 19984 13880 20036 13889
rect 20260 13923 20312 13932
rect 20260 13889 20294 13923
rect 20294 13889 20312 13923
rect 20260 13880 20312 13889
rect 20536 13880 20588 13932
rect 10232 13744 10284 13796
rect 14648 13744 14700 13796
rect 7012 13719 7064 13728
rect 7012 13685 7021 13719
rect 7021 13685 7055 13719
rect 7055 13685 7064 13719
rect 7012 13676 7064 13685
rect 9220 13676 9272 13728
rect 14556 13719 14608 13728
rect 14556 13685 14565 13719
rect 14565 13685 14599 13719
rect 14599 13685 14608 13719
rect 14556 13676 14608 13685
rect 15476 13676 15528 13728
rect 15660 13719 15712 13728
rect 15660 13685 15669 13719
rect 15669 13685 15703 13719
rect 15703 13685 15712 13719
rect 15660 13676 15712 13685
rect 17592 13787 17644 13796
rect 17592 13753 17601 13787
rect 17601 13753 17635 13787
rect 17635 13753 17644 13787
rect 17592 13744 17644 13753
rect 21364 13719 21416 13728
rect 21364 13685 21373 13719
rect 21373 13685 21407 13719
rect 21407 13685 21416 13719
rect 21364 13676 21416 13685
rect 3595 13574 3647 13626
rect 3659 13574 3711 13626
rect 3723 13574 3775 13626
rect 3787 13574 3839 13626
rect 3851 13574 3903 13626
rect 8885 13574 8937 13626
rect 8949 13574 9001 13626
rect 9013 13574 9065 13626
rect 9077 13574 9129 13626
rect 9141 13574 9193 13626
rect 14175 13574 14227 13626
rect 14239 13574 14291 13626
rect 14303 13574 14355 13626
rect 14367 13574 14419 13626
rect 14431 13574 14483 13626
rect 19465 13574 19517 13626
rect 19529 13574 19581 13626
rect 19593 13574 19645 13626
rect 19657 13574 19709 13626
rect 19721 13574 19773 13626
rect 7104 13472 7156 13524
rect 9404 13515 9456 13524
rect 9404 13481 9413 13515
rect 9413 13481 9447 13515
rect 9447 13481 9456 13515
rect 9404 13472 9456 13481
rect 9312 13447 9364 13456
rect 9312 13413 9321 13447
rect 9321 13413 9355 13447
rect 9355 13413 9364 13447
rect 9312 13404 9364 13413
rect 15476 13472 15528 13524
rect 15568 13472 15620 13524
rect 15660 13515 15712 13524
rect 15660 13481 15669 13515
rect 15669 13481 15703 13515
rect 15703 13481 15712 13515
rect 15660 13472 15712 13481
rect 4344 13336 4396 13388
rect 9220 13336 9272 13388
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 10508 13336 10560 13388
rect 12072 13336 12124 13388
rect 6000 13268 6052 13320
rect 7840 13311 7892 13320
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 10140 13268 10192 13320
rect 7472 13200 7524 13252
rect 6920 13132 6972 13184
rect 10784 13200 10836 13252
rect 11980 13200 12032 13252
rect 17592 13268 17644 13320
rect 18696 13311 18748 13320
rect 18696 13277 18705 13311
rect 18705 13277 18739 13311
rect 18739 13277 18748 13311
rect 18696 13268 18748 13277
rect 16488 13200 16540 13252
rect 18052 13200 18104 13252
rect 20628 13268 20680 13320
rect 20720 13311 20772 13320
rect 20720 13277 20729 13311
rect 20729 13277 20763 13311
rect 20763 13277 20772 13311
rect 20720 13268 20772 13277
rect 21364 13268 21416 13320
rect 13820 13132 13872 13184
rect 14556 13132 14608 13184
rect 15384 13132 15436 13184
rect 19248 13175 19300 13184
rect 19248 13141 19257 13175
rect 19257 13141 19291 13175
rect 19291 13141 19300 13175
rect 19248 13132 19300 13141
rect 19708 13175 19760 13184
rect 19708 13141 19717 13175
rect 19717 13141 19751 13175
rect 19751 13141 19760 13175
rect 19708 13132 19760 13141
rect 19800 13175 19852 13184
rect 19800 13141 19809 13175
rect 19809 13141 19843 13175
rect 19843 13141 19852 13175
rect 19800 13132 19852 13141
rect 4255 13030 4307 13082
rect 4319 13030 4371 13082
rect 4383 13030 4435 13082
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 9545 13030 9597 13082
rect 9609 13030 9661 13082
rect 9673 13030 9725 13082
rect 9737 13030 9789 13082
rect 9801 13030 9853 13082
rect 14835 13030 14887 13082
rect 14899 13030 14951 13082
rect 14963 13030 15015 13082
rect 15027 13030 15079 13082
rect 15091 13030 15143 13082
rect 20125 13030 20177 13082
rect 20189 13030 20241 13082
rect 20253 13030 20305 13082
rect 20317 13030 20369 13082
rect 20381 13030 20433 13082
rect 7012 12928 7064 12980
rect 7380 12928 7432 12980
rect 11796 12928 11848 12980
rect 6828 12903 6880 12912
rect 6828 12869 6837 12903
rect 6837 12869 6871 12903
rect 6871 12869 6880 12903
rect 6828 12860 6880 12869
rect 3516 12767 3568 12776
rect 3516 12733 3525 12767
rect 3525 12733 3559 12767
rect 3559 12733 3568 12767
rect 3516 12724 3568 12733
rect 2872 12656 2924 12708
rect 6920 12792 6972 12844
rect 7104 12835 7156 12844
rect 7104 12801 7113 12835
rect 7113 12801 7147 12835
rect 7147 12801 7156 12835
rect 7104 12792 7156 12801
rect 11704 12903 11756 12912
rect 11704 12869 11713 12903
rect 11713 12869 11747 12903
rect 11747 12869 11756 12903
rect 11704 12860 11756 12869
rect 14556 12860 14608 12912
rect 16488 12971 16540 12980
rect 16488 12937 16497 12971
rect 16497 12937 16531 12971
rect 16531 12937 16540 12971
rect 16488 12928 16540 12937
rect 19984 12928 20036 12980
rect 20628 12928 20680 12980
rect 14740 12860 14792 12912
rect 19800 12860 19852 12912
rect 15292 12835 15344 12844
rect 4068 12656 4120 12708
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 15660 12792 15712 12844
rect 16028 12835 16080 12844
rect 16028 12801 16037 12835
rect 16037 12801 16071 12835
rect 16071 12801 16080 12835
rect 16028 12792 16080 12801
rect 15384 12767 15436 12776
rect 15384 12733 15393 12767
rect 15393 12733 15427 12767
rect 15427 12733 15436 12767
rect 15384 12724 15436 12733
rect 18052 12792 18104 12844
rect 14648 12656 14700 12708
rect 19708 12724 19760 12776
rect 4436 12588 4488 12640
rect 17500 12588 17552 12640
rect 21456 12588 21508 12640
rect 3595 12486 3647 12538
rect 3659 12486 3711 12538
rect 3723 12486 3775 12538
rect 3787 12486 3839 12538
rect 3851 12486 3903 12538
rect 8885 12486 8937 12538
rect 8949 12486 9001 12538
rect 9013 12486 9065 12538
rect 9077 12486 9129 12538
rect 9141 12486 9193 12538
rect 14175 12486 14227 12538
rect 14239 12486 14291 12538
rect 14303 12486 14355 12538
rect 14367 12486 14419 12538
rect 14431 12486 14483 12538
rect 19465 12486 19517 12538
rect 19529 12486 19581 12538
rect 19593 12486 19645 12538
rect 19657 12486 19709 12538
rect 19721 12486 19773 12538
rect 3516 12384 3568 12436
rect 5540 12384 5592 12436
rect 5816 12384 5868 12436
rect 10416 12384 10468 12436
rect 10508 12427 10560 12436
rect 10508 12393 10517 12427
rect 10517 12393 10551 12427
rect 10551 12393 10560 12427
rect 10508 12384 10560 12393
rect 11980 12427 12032 12436
rect 11980 12393 11989 12427
rect 11989 12393 12023 12427
rect 12023 12393 12032 12427
rect 11980 12384 12032 12393
rect 17592 12384 17644 12436
rect 19984 12384 20036 12436
rect 3424 12359 3476 12368
rect 3424 12325 3433 12359
rect 3433 12325 3467 12359
rect 3467 12325 3476 12359
rect 3424 12316 3476 12325
rect 4068 12316 4120 12368
rect 1584 12180 1636 12232
rect 4160 12180 4212 12232
rect 4436 12180 4488 12232
rect 5264 12223 5316 12232
rect 5264 12189 5273 12223
rect 5273 12189 5307 12223
rect 5307 12189 5316 12223
rect 5264 12180 5316 12189
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 5724 12223 5776 12232
rect 5724 12189 5733 12223
rect 5733 12189 5767 12223
rect 5767 12189 5776 12223
rect 5724 12180 5776 12189
rect 9956 12180 10008 12232
rect 13820 12248 13872 12300
rect 18696 12316 18748 12368
rect 2136 12112 2188 12164
rect 10324 12112 10376 12164
rect 4620 12044 4672 12096
rect 4896 12044 4948 12096
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 8668 12044 8720 12096
rect 14556 12180 14608 12232
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 10784 12044 10836 12096
rect 11244 12044 11296 12096
rect 11888 12044 11940 12096
rect 15936 12112 15988 12164
rect 12992 12044 13044 12096
rect 13912 12044 13964 12096
rect 14004 12044 14056 12096
rect 19892 12180 19944 12232
rect 20720 12384 20772 12436
rect 21456 12427 21508 12436
rect 21456 12393 21465 12427
rect 21465 12393 21499 12427
rect 21499 12393 21508 12427
rect 21456 12384 21508 12393
rect 19156 12044 19208 12096
rect 20720 12223 20772 12232
rect 20720 12189 20729 12223
rect 20729 12189 20763 12223
rect 20763 12189 20772 12223
rect 20720 12180 20772 12189
rect 20996 12112 21048 12164
rect 20536 12044 20588 12096
rect 4255 11942 4307 11994
rect 4319 11942 4371 11994
rect 4383 11942 4435 11994
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 9545 11942 9597 11994
rect 9609 11942 9661 11994
rect 9673 11942 9725 11994
rect 9737 11942 9789 11994
rect 9801 11942 9853 11994
rect 14835 11942 14887 11994
rect 14899 11942 14951 11994
rect 14963 11942 15015 11994
rect 15027 11942 15079 11994
rect 15091 11942 15143 11994
rect 20125 11942 20177 11994
rect 20189 11942 20241 11994
rect 20253 11942 20305 11994
rect 20317 11942 20369 11994
rect 20381 11942 20433 11994
rect 4620 11840 4672 11892
rect 5540 11883 5592 11892
rect 5540 11849 5549 11883
rect 5549 11849 5583 11883
rect 5583 11849 5592 11883
rect 5540 11840 5592 11849
rect 8668 11883 8720 11892
rect 8668 11849 8677 11883
rect 8677 11849 8711 11883
rect 8711 11849 8720 11883
rect 8668 11840 8720 11849
rect 6368 11815 6420 11824
rect 6368 11781 6377 11815
rect 6377 11781 6411 11815
rect 6411 11781 6420 11815
rect 6368 11772 6420 11781
rect 6736 11772 6788 11824
rect 9680 11840 9732 11892
rect 10232 11840 10284 11892
rect 10324 11883 10376 11892
rect 10324 11849 10333 11883
rect 10333 11849 10367 11883
rect 10367 11849 10376 11883
rect 10324 11840 10376 11849
rect 10876 11840 10928 11892
rect 12992 11840 13044 11892
rect 1584 11704 1636 11756
rect 1768 11747 1820 11756
rect 1768 11713 1802 11747
rect 1802 11713 1820 11747
rect 1768 11704 1820 11713
rect 4160 11704 4212 11756
rect 3332 11568 3384 11620
rect 6184 11679 6236 11688
rect 6184 11645 6193 11679
rect 6193 11645 6227 11679
rect 6227 11645 6236 11679
rect 6184 11636 6236 11645
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 8024 11704 8076 11756
rect 10140 11772 10192 11824
rect 9772 11636 9824 11688
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 12532 11747 12584 11756
rect 12532 11713 12541 11747
rect 12541 11713 12575 11747
rect 12575 11713 12584 11747
rect 12532 11704 12584 11713
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 3056 11500 3108 11552
rect 4252 11500 4304 11552
rect 10416 11568 10468 11620
rect 12256 11679 12308 11688
rect 12256 11645 12265 11679
rect 12265 11645 12299 11679
rect 12299 11645 12308 11679
rect 12256 11636 12308 11645
rect 12808 11568 12860 11620
rect 5908 11500 5960 11552
rect 6552 11543 6604 11552
rect 6552 11509 6561 11543
rect 6561 11509 6595 11543
rect 6595 11509 6604 11543
rect 6552 11500 6604 11509
rect 7288 11500 7340 11552
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 11796 11500 11848 11552
rect 12348 11543 12400 11552
rect 12348 11509 12357 11543
rect 12357 11509 12391 11543
rect 12391 11509 12400 11543
rect 12348 11500 12400 11509
rect 14004 11772 14056 11824
rect 15752 11840 15804 11892
rect 14648 11772 14700 11824
rect 15936 11815 15988 11824
rect 15936 11781 15945 11815
rect 15945 11781 15979 11815
rect 15979 11781 15988 11815
rect 15936 11772 15988 11781
rect 16764 11772 16816 11824
rect 19248 11772 19300 11824
rect 20536 11840 20588 11892
rect 20720 11840 20772 11892
rect 16028 11704 16080 11756
rect 17592 11704 17644 11756
rect 14372 11636 14424 11688
rect 17224 11679 17276 11688
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 19248 11636 19300 11688
rect 20996 11815 21048 11824
rect 20996 11781 21005 11815
rect 21005 11781 21039 11815
rect 21039 11781 21048 11815
rect 20996 11772 21048 11781
rect 21272 11747 21324 11756
rect 21272 11713 21281 11747
rect 21281 11713 21315 11747
rect 21315 11713 21324 11747
rect 21272 11704 21324 11713
rect 20720 11636 20772 11688
rect 22192 11636 22244 11688
rect 16488 11543 16540 11552
rect 16488 11509 16497 11543
rect 16497 11509 16531 11543
rect 16531 11509 16540 11543
rect 16488 11500 16540 11509
rect 19800 11500 19852 11552
rect 3595 11398 3647 11450
rect 3659 11398 3711 11450
rect 3723 11398 3775 11450
rect 3787 11398 3839 11450
rect 3851 11398 3903 11450
rect 8885 11398 8937 11450
rect 8949 11398 9001 11450
rect 9013 11398 9065 11450
rect 9077 11398 9129 11450
rect 9141 11398 9193 11450
rect 14175 11398 14227 11450
rect 14239 11398 14291 11450
rect 14303 11398 14355 11450
rect 14367 11398 14419 11450
rect 14431 11398 14483 11450
rect 19465 11398 19517 11450
rect 19529 11398 19581 11450
rect 19593 11398 19645 11450
rect 19657 11398 19709 11450
rect 19721 11398 19773 11450
rect 1768 11296 1820 11348
rect 2136 11339 2188 11348
rect 2136 11305 2145 11339
rect 2145 11305 2179 11339
rect 2179 11305 2188 11339
rect 2136 11296 2188 11305
rect 2872 11296 2924 11348
rect 3056 11296 3108 11348
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 4252 11296 4304 11348
rect 6552 11296 6604 11348
rect 9772 11339 9824 11348
rect 6368 11228 6420 11280
rect 6644 11228 6696 11280
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 2780 11092 2832 11144
rect 2964 10956 3016 11008
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 3516 11092 3568 11144
rect 4160 11160 4212 11212
rect 4620 11203 4672 11212
rect 4620 11169 4629 11203
rect 4629 11169 4663 11203
rect 4663 11169 4672 11203
rect 4620 11160 4672 11169
rect 6828 11160 6880 11212
rect 9772 11305 9781 11339
rect 9781 11305 9815 11339
rect 9815 11305 9824 11339
rect 9772 11296 9824 11305
rect 8760 11228 8812 11280
rect 4896 11135 4948 11144
rect 4896 11101 4930 11135
rect 4930 11101 4948 11135
rect 4896 11092 4948 11101
rect 6368 11135 6420 11144
rect 6368 11101 6377 11135
rect 6377 11101 6411 11135
rect 6411 11101 6420 11135
rect 6368 11092 6420 11101
rect 9956 11092 10008 11144
rect 10600 11296 10652 11348
rect 12624 11296 12676 11348
rect 14556 11296 14608 11348
rect 14648 11296 14700 11348
rect 13544 11160 13596 11212
rect 10968 11092 11020 11144
rect 3332 10956 3384 11008
rect 7748 11024 7800 11076
rect 9588 11024 9640 11076
rect 3884 10956 3936 11008
rect 6184 10956 6236 11008
rect 6552 10956 6604 11008
rect 7012 10999 7064 11008
rect 7012 10965 7021 10999
rect 7021 10965 7055 10999
rect 7055 10965 7064 10999
rect 7012 10956 7064 10965
rect 10140 10999 10192 11008
rect 10140 10965 10149 10999
rect 10149 10965 10183 10999
rect 10183 10965 10192 10999
rect 10140 10956 10192 10965
rect 11152 11024 11204 11076
rect 11244 11024 11296 11076
rect 12348 11024 12400 11076
rect 12256 10956 12308 11008
rect 13544 10999 13596 11008
rect 13544 10965 13553 10999
rect 13553 10965 13587 10999
rect 13587 10965 13596 10999
rect 13544 10956 13596 10965
rect 13636 10999 13688 11008
rect 13636 10965 13645 10999
rect 13645 10965 13679 10999
rect 13679 10965 13688 10999
rect 13636 10956 13688 10965
rect 14556 11024 14608 11076
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 17592 11160 17644 11212
rect 18236 11160 18288 11212
rect 19156 11296 19208 11348
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 19800 11296 19852 11348
rect 21272 11296 21324 11348
rect 21364 11296 21416 11348
rect 19340 11228 19392 11280
rect 19892 11228 19944 11280
rect 20628 11160 20680 11212
rect 15384 11024 15436 11076
rect 15660 11024 15712 11076
rect 13820 10956 13872 11008
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 16856 11024 16908 11076
rect 20536 11024 20588 11076
rect 20628 11067 20680 11076
rect 20628 11033 20653 11067
rect 20653 11033 20680 11067
rect 20628 11024 20680 11033
rect 17224 10956 17276 11008
rect 19800 10956 19852 11008
rect 4255 10854 4307 10906
rect 4319 10854 4371 10906
rect 4383 10854 4435 10906
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 9545 10854 9597 10906
rect 9609 10854 9661 10906
rect 9673 10854 9725 10906
rect 9737 10854 9789 10906
rect 9801 10854 9853 10906
rect 14835 10854 14887 10906
rect 14899 10854 14951 10906
rect 14963 10854 15015 10906
rect 15027 10854 15079 10906
rect 15091 10854 15143 10906
rect 20125 10854 20177 10906
rect 20189 10854 20241 10906
rect 20253 10854 20305 10906
rect 20317 10854 20369 10906
rect 20381 10854 20433 10906
rect 2412 10752 2464 10804
rect 2780 10752 2832 10804
rect 6368 10752 6420 10804
rect 7104 10752 7156 10804
rect 7288 10752 7340 10804
rect 7748 10795 7800 10804
rect 7748 10761 7757 10795
rect 7757 10761 7791 10795
rect 7791 10761 7800 10795
rect 7748 10752 7800 10761
rect 8024 10795 8076 10804
rect 8024 10761 8033 10795
rect 8033 10761 8067 10795
rect 8067 10761 8076 10795
rect 8024 10752 8076 10761
rect 10140 10752 10192 10804
rect 6000 10684 6052 10736
rect 11336 10752 11388 10804
rect 12808 10795 12860 10804
rect 12808 10761 12817 10795
rect 12817 10761 12851 10795
rect 12851 10761 12860 10795
rect 12808 10752 12860 10761
rect 14556 10752 14608 10804
rect 15936 10752 15988 10804
rect 16488 10752 16540 10804
rect 3332 10616 3384 10668
rect 3884 10659 3936 10668
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 4620 10616 4672 10668
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 7012 10616 7064 10668
rect 11612 10684 11664 10736
rect 2964 10548 3016 10600
rect 5908 10548 5960 10600
rect 6828 10480 6880 10532
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 14832 10616 14884 10668
rect 15384 10616 15436 10668
rect 15660 10727 15712 10736
rect 15660 10693 15669 10727
rect 15669 10693 15703 10727
rect 15703 10693 15712 10727
rect 15660 10684 15712 10693
rect 9956 10591 10008 10600
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 9956 10548 10008 10557
rect 13452 10591 13504 10600
rect 13452 10557 13461 10591
rect 13461 10557 13495 10591
rect 13495 10557 13504 10591
rect 13452 10548 13504 10557
rect 13636 10548 13688 10600
rect 15936 10659 15988 10668
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 15936 10616 15988 10625
rect 17224 10752 17276 10804
rect 19340 10684 19392 10736
rect 16672 10659 16724 10668
rect 16672 10625 16681 10659
rect 16681 10625 16715 10659
rect 16715 10625 16724 10659
rect 16672 10616 16724 10625
rect 18236 10616 18288 10668
rect 16488 10548 16540 10600
rect 12256 10480 12308 10532
rect 1952 10412 2004 10464
rect 5724 10412 5776 10464
rect 6644 10455 6696 10464
rect 6644 10421 6653 10455
rect 6653 10421 6687 10455
rect 6687 10421 6696 10455
rect 6644 10412 6696 10421
rect 12072 10455 12124 10464
rect 12072 10421 12081 10455
rect 12081 10421 12115 10455
rect 12115 10421 12124 10455
rect 12072 10412 12124 10421
rect 15292 10412 15344 10464
rect 15752 10455 15804 10464
rect 15752 10421 15761 10455
rect 15761 10421 15795 10455
rect 15795 10421 15804 10455
rect 15752 10412 15804 10421
rect 16856 10412 16908 10464
rect 20996 10412 21048 10464
rect 21640 10455 21692 10464
rect 21640 10421 21649 10455
rect 21649 10421 21683 10455
rect 21683 10421 21692 10455
rect 21640 10412 21692 10421
rect 3595 10310 3647 10362
rect 3659 10310 3711 10362
rect 3723 10310 3775 10362
rect 3787 10310 3839 10362
rect 3851 10310 3903 10362
rect 8885 10310 8937 10362
rect 8949 10310 9001 10362
rect 9013 10310 9065 10362
rect 9077 10310 9129 10362
rect 9141 10310 9193 10362
rect 14175 10310 14227 10362
rect 14239 10310 14291 10362
rect 14303 10310 14355 10362
rect 14367 10310 14419 10362
rect 14431 10310 14483 10362
rect 19465 10310 19517 10362
rect 19529 10310 19581 10362
rect 19593 10310 19645 10362
rect 19657 10310 19709 10362
rect 19721 10310 19773 10362
rect 3332 10208 3384 10260
rect 5264 10208 5316 10260
rect 1584 10072 1636 10124
rect 5908 10072 5960 10124
rect 6736 10251 6788 10260
rect 6736 10217 6745 10251
rect 6745 10217 6779 10251
rect 6779 10217 6788 10251
rect 6736 10208 6788 10217
rect 12072 10208 12124 10260
rect 12532 10251 12584 10260
rect 12532 10217 12541 10251
rect 12541 10217 12575 10251
rect 12575 10217 12584 10251
rect 12532 10208 12584 10217
rect 12900 10208 12952 10260
rect 13636 10208 13688 10260
rect 14832 10251 14884 10260
rect 14832 10217 14841 10251
rect 14841 10217 14875 10251
rect 14875 10217 14884 10251
rect 14832 10208 14884 10217
rect 1952 10004 2004 10056
rect 5724 10004 5776 10056
rect 6368 9979 6420 9988
rect 6368 9945 6377 9979
rect 6377 9945 6411 9979
rect 6411 9945 6420 9979
rect 6368 9936 6420 9945
rect 6552 9979 6604 9988
rect 6552 9945 6577 9979
rect 6577 9945 6604 9979
rect 10048 10004 10100 10056
rect 10324 10004 10376 10056
rect 11612 10004 11664 10056
rect 12348 10047 12400 10056
rect 12348 10013 12357 10047
rect 12357 10013 12391 10047
rect 12391 10013 12400 10047
rect 12348 10004 12400 10013
rect 12624 10004 12676 10056
rect 13544 10004 13596 10056
rect 14372 10004 14424 10056
rect 15752 10208 15804 10260
rect 20536 10208 20588 10260
rect 16488 10140 16540 10192
rect 20720 10251 20772 10260
rect 20720 10217 20729 10251
rect 20729 10217 20763 10251
rect 20763 10217 20772 10251
rect 20720 10208 20772 10217
rect 21640 10208 21692 10260
rect 15384 10004 15436 10056
rect 19064 10047 19116 10056
rect 19064 10013 19073 10047
rect 19073 10013 19107 10047
rect 19107 10013 19116 10047
rect 19064 10004 19116 10013
rect 20536 10004 20588 10056
rect 20720 10004 20772 10056
rect 20904 10047 20956 10056
rect 20904 10013 20913 10047
rect 20913 10013 20947 10047
rect 20947 10013 20956 10047
rect 20904 10004 20956 10013
rect 20996 10047 21048 10056
rect 20996 10013 21005 10047
rect 21005 10013 21039 10047
rect 21039 10013 21048 10047
rect 20996 10004 21048 10013
rect 6552 9936 6604 9945
rect 12256 9936 12308 9988
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 19340 9936 19392 9988
rect 21088 9936 21140 9988
rect 17224 9868 17276 9920
rect 18420 9911 18472 9920
rect 18420 9877 18429 9911
rect 18429 9877 18463 9911
rect 18463 9877 18472 9911
rect 18420 9868 18472 9877
rect 21272 9911 21324 9920
rect 21272 9877 21281 9911
rect 21281 9877 21315 9911
rect 21315 9877 21324 9911
rect 21272 9868 21324 9877
rect 4255 9766 4307 9818
rect 4319 9766 4371 9818
rect 4383 9766 4435 9818
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 9545 9766 9597 9818
rect 9609 9766 9661 9818
rect 9673 9766 9725 9818
rect 9737 9766 9789 9818
rect 9801 9766 9853 9818
rect 14835 9766 14887 9818
rect 14899 9766 14951 9818
rect 14963 9766 15015 9818
rect 15027 9766 15079 9818
rect 15091 9766 15143 9818
rect 20125 9766 20177 9818
rect 20189 9766 20241 9818
rect 20253 9766 20305 9818
rect 20317 9766 20369 9818
rect 20381 9766 20433 9818
rect 2964 9707 3016 9716
rect 2964 9673 2973 9707
rect 2973 9673 3007 9707
rect 3007 9673 3016 9707
rect 2964 9664 3016 9673
rect 3148 9596 3200 9648
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 2228 9528 2280 9580
rect 4068 9596 4120 9648
rect 10048 9664 10100 9716
rect 12348 9664 12400 9716
rect 5540 9528 5592 9580
rect 4344 9460 4396 9512
rect 6368 9528 6420 9580
rect 7748 9528 7800 9580
rect 8300 9571 8352 9580
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 9312 9596 9364 9648
rect 10784 9596 10836 9648
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 8668 9460 8720 9512
rect 7288 9392 7340 9444
rect 3976 9367 4028 9376
rect 3976 9333 3985 9367
rect 3985 9333 4019 9367
rect 4019 9333 4028 9367
rect 3976 9324 4028 9333
rect 5080 9324 5132 9376
rect 5264 9367 5316 9376
rect 5264 9333 5273 9367
rect 5273 9333 5307 9367
rect 5307 9333 5316 9367
rect 5264 9324 5316 9333
rect 5632 9367 5684 9376
rect 5632 9333 5641 9367
rect 5641 9333 5675 9367
rect 5675 9333 5684 9367
rect 5632 9324 5684 9333
rect 6092 9367 6144 9376
rect 6092 9333 6101 9367
rect 6101 9333 6135 9367
rect 6135 9333 6144 9367
rect 6092 9324 6144 9333
rect 7380 9324 7432 9376
rect 8116 9324 8168 9376
rect 8208 9324 8260 9376
rect 8392 9367 8444 9376
rect 8392 9333 8401 9367
rect 8401 9333 8435 9367
rect 8435 9333 8444 9367
rect 8392 9324 8444 9333
rect 9956 9460 10008 9512
rect 10048 9503 10100 9512
rect 10048 9469 10058 9503
rect 10058 9469 10092 9503
rect 10092 9469 10100 9503
rect 10048 9460 10100 9469
rect 10232 9503 10284 9512
rect 10232 9469 10241 9503
rect 10241 9469 10275 9503
rect 10275 9469 10284 9503
rect 10232 9460 10284 9469
rect 10416 9528 10468 9580
rect 10600 9528 10652 9580
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 16028 9664 16080 9716
rect 14372 9596 14424 9648
rect 14556 9596 14608 9648
rect 14096 9528 14148 9580
rect 16672 9664 16724 9716
rect 19064 9664 19116 9716
rect 21088 9664 21140 9716
rect 21272 9664 21324 9716
rect 20904 9596 20956 9648
rect 18420 9571 18472 9580
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 18604 9571 18656 9580
rect 18604 9537 18613 9571
rect 18613 9537 18647 9571
rect 18647 9537 18656 9571
rect 18604 9528 18656 9537
rect 20444 9528 20496 9580
rect 10416 9392 10468 9444
rect 11888 9460 11940 9512
rect 17224 9460 17276 9512
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 19340 9392 19392 9444
rect 20628 9435 20680 9444
rect 20628 9401 20637 9435
rect 20637 9401 20671 9435
rect 20671 9401 20680 9435
rect 20628 9392 20680 9401
rect 11612 9324 11664 9376
rect 20996 9324 21048 9376
rect 21088 9367 21140 9376
rect 21088 9333 21097 9367
rect 21097 9333 21131 9367
rect 21131 9333 21140 9367
rect 21088 9324 21140 9333
rect 3595 9222 3647 9274
rect 3659 9222 3711 9274
rect 3723 9222 3775 9274
rect 3787 9222 3839 9274
rect 3851 9222 3903 9274
rect 8885 9222 8937 9274
rect 8949 9222 9001 9274
rect 9013 9222 9065 9274
rect 9077 9222 9129 9274
rect 9141 9222 9193 9274
rect 14175 9222 14227 9274
rect 14239 9222 14291 9274
rect 14303 9222 14355 9274
rect 14367 9222 14419 9274
rect 14431 9222 14483 9274
rect 19465 9222 19517 9274
rect 19529 9222 19581 9274
rect 19593 9222 19645 9274
rect 19657 9222 19709 9274
rect 19721 9222 19773 9274
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 4068 9120 4120 9172
rect 4344 9163 4396 9172
rect 4344 9129 4353 9163
rect 4353 9129 4387 9163
rect 4387 9129 4396 9163
rect 4344 9120 4396 9129
rect 5632 9120 5684 9172
rect 6092 9120 6144 9172
rect 8116 9120 8168 9172
rect 8300 9120 8352 9172
rect 940 8916 992 8968
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 4068 8916 4120 8968
rect 5540 8984 5592 9036
rect 5080 8916 5132 8968
rect 6092 8916 6144 8968
rect 8208 8916 8260 8968
rect 9036 8984 9088 9036
rect 10048 9120 10100 9172
rect 10416 9120 10468 9172
rect 11428 9120 11480 9172
rect 4160 8780 4212 8832
rect 7288 8780 7340 8832
rect 8024 8780 8076 8832
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 10508 9052 10560 9104
rect 11152 9052 11204 9104
rect 11796 9163 11848 9172
rect 11796 9129 11805 9163
rect 11805 9129 11839 9163
rect 11839 9129 11848 9163
rect 11796 9120 11848 9129
rect 11888 9163 11940 9172
rect 11888 9129 11897 9163
rect 11897 9129 11931 9163
rect 11931 9129 11940 9163
rect 11888 9120 11940 9129
rect 13544 9120 13596 9172
rect 20444 9163 20496 9172
rect 20444 9129 20453 9163
rect 20453 9129 20487 9163
rect 20487 9129 20496 9163
rect 20444 9120 20496 9129
rect 21180 9120 21232 9172
rect 10416 8984 10468 9036
rect 10232 8916 10284 8968
rect 10508 8916 10560 8968
rect 11244 8984 11296 9036
rect 11336 9027 11388 9036
rect 11336 8993 11345 9027
rect 11345 8993 11379 9027
rect 11379 8993 11388 9027
rect 11336 8984 11388 8993
rect 11428 9027 11480 9036
rect 11428 8993 11437 9027
rect 11437 8993 11471 9027
rect 11471 8993 11480 9027
rect 11428 8984 11480 8993
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 11704 8916 11756 8968
rect 12072 8959 12124 8968
rect 12072 8925 12081 8959
rect 12081 8925 12115 8959
rect 12115 8925 12124 8959
rect 12072 8916 12124 8925
rect 9496 8848 9548 8900
rect 8668 8780 8720 8832
rect 9128 8780 9180 8832
rect 9312 8780 9364 8832
rect 12716 8916 12768 8968
rect 19984 9052 20036 9104
rect 10140 8823 10192 8832
rect 10140 8789 10149 8823
rect 10149 8789 10183 8823
rect 10183 8789 10192 8823
rect 10140 8780 10192 8789
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 11060 8780 11112 8832
rect 15384 8916 15436 8968
rect 16120 8916 16172 8968
rect 16856 8916 16908 8968
rect 20536 9027 20588 9036
rect 20536 8993 20545 9027
rect 20545 8993 20579 9027
rect 20579 8993 20588 9027
rect 20536 8984 20588 8993
rect 17408 8959 17460 8968
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 15200 8891 15252 8900
rect 15200 8857 15218 8891
rect 15218 8857 15252 8891
rect 15200 8848 15252 8857
rect 21088 8916 21140 8968
rect 20720 8848 20772 8900
rect 12348 8780 12400 8832
rect 13452 8780 13504 8832
rect 16580 8780 16632 8832
rect 4255 8678 4307 8730
rect 4319 8678 4371 8730
rect 4383 8678 4435 8730
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 9545 8678 9597 8730
rect 9609 8678 9661 8730
rect 9673 8678 9725 8730
rect 9737 8678 9789 8730
rect 9801 8678 9853 8730
rect 14835 8678 14887 8730
rect 14899 8678 14951 8730
rect 14963 8678 15015 8730
rect 15027 8678 15079 8730
rect 15091 8678 15143 8730
rect 20125 8678 20177 8730
rect 20189 8678 20241 8730
rect 20253 8678 20305 8730
rect 20317 8678 20369 8730
rect 20381 8678 20433 8730
rect 3976 8576 4028 8628
rect 5264 8576 5316 8628
rect 6092 8619 6144 8628
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 9036 8576 9088 8628
rect 9404 8576 9456 8628
rect 9956 8576 10008 8628
rect 10600 8576 10652 8628
rect 10692 8576 10744 8628
rect 11336 8619 11388 8628
rect 11336 8585 11345 8619
rect 11345 8585 11379 8619
rect 11379 8585 11388 8619
rect 11336 8576 11388 8585
rect 7012 8508 7064 8560
rect 1584 8440 1636 8492
rect 7380 8440 7432 8492
rect 7656 8440 7708 8492
rect 8300 8483 8352 8492
rect 8300 8449 8309 8483
rect 8309 8449 8343 8483
rect 8343 8449 8352 8483
rect 8300 8440 8352 8449
rect 9128 8551 9180 8560
rect 9128 8517 9137 8551
rect 9137 8517 9171 8551
rect 9171 8517 9180 8551
rect 9128 8508 9180 8517
rect 6920 8415 6972 8424
rect 6920 8381 6929 8415
rect 6929 8381 6963 8415
rect 6963 8381 6972 8415
rect 6920 8372 6972 8381
rect 7840 8372 7892 8424
rect 8668 8372 8720 8424
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 9864 8508 9916 8560
rect 9588 8440 9640 8492
rect 3516 8236 3568 8288
rect 8392 8304 8444 8356
rect 8484 8347 8536 8356
rect 8484 8313 8493 8347
rect 8493 8313 8527 8347
rect 8527 8313 8536 8347
rect 8484 8304 8536 8313
rect 9404 8304 9456 8356
rect 5080 8236 5132 8288
rect 9312 8236 9364 8288
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 11704 8576 11756 8628
rect 12716 8576 12768 8628
rect 10692 8372 10744 8424
rect 11428 8372 11480 8424
rect 11612 8440 11664 8492
rect 13636 8483 13688 8492
rect 13636 8449 13645 8483
rect 13645 8449 13679 8483
rect 13679 8449 13688 8483
rect 13636 8440 13688 8449
rect 16120 8576 16172 8628
rect 15384 8508 15436 8560
rect 17408 8576 17460 8628
rect 19892 8576 19944 8628
rect 14096 8440 14148 8492
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 16580 8440 16632 8492
rect 21180 8440 21232 8492
rect 9588 8304 9640 8356
rect 11060 8304 11112 8356
rect 10232 8279 10284 8288
rect 10232 8245 10241 8279
rect 10241 8245 10275 8279
rect 10275 8245 10284 8279
rect 10232 8236 10284 8245
rect 10416 8236 10468 8288
rect 10968 8236 11020 8288
rect 13452 8347 13504 8356
rect 13452 8313 13461 8347
rect 13461 8313 13495 8347
rect 13495 8313 13504 8347
rect 13452 8304 13504 8313
rect 17684 8372 17736 8424
rect 13728 8236 13780 8288
rect 13820 8279 13872 8288
rect 13820 8245 13829 8279
rect 13829 8245 13863 8279
rect 13863 8245 13872 8279
rect 13820 8236 13872 8245
rect 15292 8236 15344 8288
rect 15476 8236 15528 8288
rect 16396 8236 16448 8288
rect 18052 8279 18104 8288
rect 18052 8245 18061 8279
rect 18061 8245 18095 8279
rect 18095 8245 18104 8279
rect 18052 8236 18104 8245
rect 18604 8236 18656 8288
rect 3595 8134 3647 8186
rect 3659 8134 3711 8186
rect 3723 8134 3775 8186
rect 3787 8134 3839 8186
rect 3851 8134 3903 8186
rect 8885 8134 8937 8186
rect 8949 8134 9001 8186
rect 9013 8134 9065 8186
rect 9077 8134 9129 8186
rect 9141 8134 9193 8186
rect 14175 8134 14227 8186
rect 14239 8134 14291 8186
rect 14303 8134 14355 8186
rect 14367 8134 14419 8186
rect 14431 8134 14483 8186
rect 19465 8134 19517 8186
rect 19529 8134 19581 8186
rect 19593 8134 19645 8186
rect 19657 8134 19709 8186
rect 19721 8134 19773 8186
rect 6092 7964 6144 8016
rect 3516 7828 3568 7880
rect 3884 7828 3936 7880
rect 4160 7760 4212 7812
rect 6920 7896 6972 7948
rect 7472 7964 7524 8016
rect 5356 7828 5408 7880
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 7656 8075 7708 8084
rect 7656 8041 7665 8075
rect 7665 8041 7699 8075
rect 7699 8041 7708 8075
rect 7656 8032 7708 8041
rect 7748 8032 7800 8084
rect 9220 8032 9272 8084
rect 10324 8032 10376 8084
rect 11428 8032 11480 8084
rect 7840 7896 7892 7948
rect 8024 7896 8076 7948
rect 9588 7964 9640 8016
rect 12072 8075 12124 8084
rect 12072 8041 12081 8075
rect 12081 8041 12115 8075
rect 12115 8041 12124 8075
rect 12072 8032 12124 8041
rect 13636 8032 13688 8084
rect 14096 8032 14148 8084
rect 14556 8032 14608 8084
rect 15200 8032 15252 8084
rect 13820 7964 13872 8016
rect 9956 7896 10008 7948
rect 10324 7896 10376 7948
rect 6828 7760 6880 7812
rect 8024 7803 8076 7812
rect 8024 7769 8043 7803
rect 8043 7769 8076 7803
rect 10048 7828 10100 7880
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 10232 7828 10284 7880
rect 10416 7828 10468 7880
rect 12348 7871 12400 7880
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 12440 7871 12492 7880
rect 12440 7837 12449 7871
rect 12449 7837 12483 7871
rect 12483 7837 12492 7871
rect 12440 7828 12492 7837
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 12624 7871 12676 7880
rect 12624 7837 12633 7871
rect 12633 7837 12667 7871
rect 12667 7837 12676 7871
rect 12624 7828 12676 7837
rect 17684 8075 17736 8084
rect 17684 8041 17693 8075
rect 17693 8041 17727 8075
rect 17727 8041 17736 8075
rect 17684 8032 17736 8041
rect 18972 7964 19024 8016
rect 15384 7896 15436 7948
rect 18052 7939 18104 7948
rect 18052 7905 18061 7939
rect 18061 7905 18095 7939
rect 18095 7905 18104 7939
rect 18052 7896 18104 7905
rect 8024 7760 8076 7769
rect 5172 7735 5224 7744
rect 5172 7701 5181 7735
rect 5181 7701 5215 7735
rect 5215 7701 5224 7735
rect 5172 7692 5224 7701
rect 5540 7692 5592 7744
rect 6920 7692 6972 7744
rect 8760 7692 8812 7744
rect 9864 7692 9916 7744
rect 11980 7760 12032 7812
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 19340 7828 19392 7880
rect 14556 7692 14608 7744
rect 16672 7760 16724 7812
rect 20628 7828 20680 7880
rect 20720 7828 20772 7880
rect 21824 7871 21876 7880
rect 21824 7837 21833 7871
rect 21833 7837 21867 7871
rect 21867 7837 21876 7871
rect 21824 7828 21876 7837
rect 18420 7692 18472 7744
rect 19248 7735 19300 7744
rect 19248 7701 19257 7735
rect 19257 7701 19291 7735
rect 19291 7701 19300 7735
rect 19248 7692 19300 7701
rect 20812 7692 20864 7744
rect 21548 7692 21600 7744
rect 4255 7590 4307 7642
rect 4319 7590 4371 7642
rect 4383 7590 4435 7642
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 9545 7590 9597 7642
rect 9609 7590 9661 7642
rect 9673 7590 9725 7642
rect 9737 7590 9789 7642
rect 9801 7590 9853 7642
rect 14835 7590 14887 7642
rect 14899 7590 14951 7642
rect 14963 7590 15015 7642
rect 15027 7590 15079 7642
rect 15091 7590 15143 7642
rect 20125 7590 20177 7642
rect 20189 7590 20241 7642
rect 20253 7590 20305 7642
rect 20317 7590 20369 7642
rect 20381 7590 20433 7642
rect 5080 7488 5132 7540
rect 5264 7420 5316 7472
rect 6092 7488 6144 7540
rect 7012 7488 7064 7540
rect 7104 7488 7156 7540
rect 5172 7352 5224 7404
rect 3976 7148 4028 7200
rect 6828 7420 6880 7472
rect 11704 7488 11756 7540
rect 11980 7488 12032 7540
rect 12440 7488 12492 7540
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 8392 7352 8444 7404
rect 14556 7463 14608 7472
rect 13912 7352 13964 7404
rect 14556 7429 14565 7463
rect 14565 7429 14599 7463
rect 14599 7429 14608 7463
rect 14556 7420 14608 7429
rect 14648 7352 14700 7404
rect 5724 7191 5776 7200
rect 5724 7157 5733 7191
rect 5733 7157 5767 7191
rect 5767 7157 5776 7191
rect 5724 7148 5776 7157
rect 8300 7284 8352 7336
rect 12072 7284 12124 7336
rect 15292 7284 15344 7336
rect 17500 7327 17552 7336
rect 17500 7293 17509 7327
rect 17509 7293 17543 7327
rect 17543 7293 17552 7327
rect 17500 7284 17552 7293
rect 18052 7284 18104 7336
rect 10324 7148 10376 7200
rect 12624 7148 12676 7200
rect 16948 7148 17000 7200
rect 19248 7352 19300 7404
rect 19984 7420 20036 7472
rect 20628 7488 20680 7540
rect 20536 7420 20588 7472
rect 20168 7352 20220 7404
rect 20628 7352 20680 7404
rect 21548 7352 21600 7404
rect 19892 7327 19944 7336
rect 19892 7293 19901 7327
rect 19901 7293 19935 7327
rect 19935 7293 19944 7327
rect 19892 7284 19944 7293
rect 20444 7148 20496 7200
rect 3595 7046 3647 7098
rect 3659 7046 3711 7098
rect 3723 7046 3775 7098
rect 3787 7046 3839 7098
rect 3851 7046 3903 7098
rect 8885 7046 8937 7098
rect 8949 7046 9001 7098
rect 9013 7046 9065 7098
rect 9077 7046 9129 7098
rect 9141 7046 9193 7098
rect 14175 7046 14227 7098
rect 14239 7046 14291 7098
rect 14303 7046 14355 7098
rect 14367 7046 14419 7098
rect 14431 7046 14483 7098
rect 19465 7046 19517 7098
rect 19529 7046 19581 7098
rect 19593 7046 19645 7098
rect 19657 7046 19709 7098
rect 19721 7046 19773 7098
rect 8024 6944 8076 6996
rect 4068 6740 4120 6792
rect 7196 6808 7248 6860
rect 8484 6808 8536 6860
rect 7288 6740 7340 6792
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 8576 6740 8628 6792
rect 9864 6808 9916 6860
rect 5724 6672 5776 6724
rect 6460 6672 6512 6724
rect 8208 6715 8260 6724
rect 8208 6681 8217 6715
rect 8217 6681 8251 6715
rect 8251 6681 8260 6715
rect 8208 6672 8260 6681
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 9404 6740 9456 6792
rect 9864 6715 9916 6724
rect 9864 6681 9873 6715
rect 9873 6681 9907 6715
rect 9907 6681 9916 6715
rect 9864 6672 9916 6681
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 4896 6647 4948 6656
rect 4896 6613 4905 6647
rect 4905 6613 4939 6647
rect 4939 6613 4948 6647
rect 4896 6604 4948 6613
rect 8392 6604 8444 6656
rect 8668 6604 8720 6656
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 12532 6944 12584 6996
rect 16672 6987 16724 6996
rect 16672 6953 16681 6987
rect 16681 6953 16715 6987
rect 16715 6953 16724 6987
rect 16672 6944 16724 6953
rect 17592 6944 17644 6996
rect 17960 6987 18012 6996
rect 17960 6953 17969 6987
rect 17969 6953 18003 6987
rect 18003 6953 18012 6987
rect 17960 6944 18012 6953
rect 18052 6944 18104 6996
rect 19340 6944 19392 6996
rect 11152 6808 11204 6860
rect 17684 6919 17736 6928
rect 17684 6885 17693 6919
rect 17693 6885 17727 6919
rect 17727 6885 17736 6919
rect 17684 6876 17736 6885
rect 13912 6808 13964 6860
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 12072 6740 12124 6792
rect 14556 6740 14608 6792
rect 16120 6808 16172 6860
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 19892 6987 19944 6996
rect 19892 6953 19901 6987
rect 19901 6953 19935 6987
rect 19935 6953 19944 6987
rect 19892 6944 19944 6953
rect 20536 6851 20588 6860
rect 20536 6817 20545 6851
rect 20545 6817 20579 6851
rect 20579 6817 20588 6851
rect 20536 6808 20588 6817
rect 15844 6740 15896 6792
rect 16856 6783 16908 6792
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 16856 6740 16908 6749
rect 16948 6783 17000 6792
rect 16948 6749 16957 6783
rect 16957 6749 16991 6783
rect 16991 6749 17000 6783
rect 16948 6740 17000 6749
rect 17500 6740 17552 6792
rect 10048 6604 10100 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 14648 6604 14700 6656
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 16856 6604 16908 6656
rect 17408 6647 17460 6656
rect 17408 6613 17417 6647
rect 17417 6613 17451 6647
rect 17451 6613 17460 6647
rect 17408 6604 17460 6613
rect 17592 6672 17644 6724
rect 17684 6672 17736 6724
rect 17868 6672 17920 6724
rect 18420 6783 18472 6792
rect 18420 6749 18429 6783
rect 18429 6749 18463 6783
rect 18463 6749 18472 6783
rect 18420 6740 18472 6749
rect 20812 6783 20864 6792
rect 19984 6672 20036 6724
rect 20812 6749 20846 6783
rect 20846 6749 20864 6783
rect 20812 6740 20864 6749
rect 18052 6604 18104 6656
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 18788 6604 18840 6613
rect 20168 6604 20220 6656
rect 20444 6604 20496 6656
rect 4255 6502 4307 6554
rect 4319 6502 4371 6554
rect 4383 6502 4435 6554
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 9545 6502 9597 6554
rect 9609 6502 9661 6554
rect 9673 6502 9725 6554
rect 9737 6502 9789 6554
rect 9801 6502 9853 6554
rect 14835 6502 14887 6554
rect 14899 6502 14951 6554
rect 14963 6502 15015 6554
rect 15027 6502 15079 6554
rect 15091 6502 15143 6554
rect 20125 6502 20177 6554
rect 20189 6502 20241 6554
rect 20253 6502 20305 6554
rect 20317 6502 20369 6554
rect 20381 6502 20433 6554
rect 4068 6400 4120 6452
rect 4160 6400 4212 6452
rect 4896 6332 4948 6384
rect 7196 6400 7248 6452
rect 7288 6400 7340 6452
rect 8392 6400 8444 6452
rect 8576 6400 8628 6452
rect 9220 6443 9272 6452
rect 9220 6409 9229 6443
rect 9229 6409 9263 6443
rect 9263 6409 9272 6443
rect 9220 6400 9272 6409
rect 10048 6400 10100 6452
rect 10416 6400 10468 6452
rect 11520 6400 11572 6452
rect 11888 6400 11940 6452
rect 8024 6332 8076 6384
rect 3240 6196 3292 6248
rect 5540 6239 5592 6248
rect 5540 6205 5549 6239
rect 5549 6205 5583 6239
rect 5583 6205 5592 6239
rect 5540 6196 5592 6205
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 6920 6196 6972 6205
rect 7104 6307 7156 6316
rect 7104 6273 7113 6307
rect 7113 6273 7147 6307
rect 7147 6273 7156 6307
rect 7104 6264 7156 6273
rect 7564 6264 7616 6316
rect 7380 6196 7432 6248
rect 7840 6239 7892 6248
rect 7840 6205 7849 6239
rect 7849 6205 7883 6239
rect 7883 6205 7892 6239
rect 7840 6196 7892 6205
rect 7380 6060 7432 6112
rect 8208 6196 8260 6248
rect 8760 6264 8812 6316
rect 9312 6264 9364 6316
rect 13912 6443 13964 6452
rect 13912 6409 13921 6443
rect 13921 6409 13955 6443
rect 13955 6409 13964 6443
rect 13912 6400 13964 6409
rect 14096 6400 14148 6452
rect 12624 6375 12676 6384
rect 12624 6341 12633 6375
rect 12633 6341 12667 6375
rect 12667 6341 12676 6375
rect 12624 6332 12676 6341
rect 13268 6332 13320 6384
rect 15476 6400 15528 6452
rect 12072 6264 12124 6316
rect 9220 6196 9272 6248
rect 9588 6239 9640 6248
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 9864 6196 9916 6248
rect 8300 6128 8352 6180
rect 9588 6060 9640 6112
rect 12164 6128 12216 6180
rect 15292 6239 15344 6248
rect 15292 6205 15301 6239
rect 15301 6205 15335 6239
rect 15335 6205 15344 6239
rect 15292 6196 15344 6205
rect 17408 6400 17460 6452
rect 17776 6400 17828 6452
rect 17868 6400 17920 6452
rect 19892 6400 19944 6452
rect 13268 6171 13320 6180
rect 13268 6137 13277 6171
rect 13277 6137 13311 6171
rect 13311 6137 13320 6171
rect 13268 6128 13320 6137
rect 16028 6196 16080 6248
rect 17868 6264 17920 6316
rect 18788 6264 18840 6316
rect 19984 6332 20036 6384
rect 20536 6332 20588 6384
rect 20260 6264 20312 6316
rect 11152 6060 11204 6112
rect 13084 6103 13136 6112
rect 13084 6069 13093 6103
rect 13093 6069 13127 6103
rect 13127 6069 13136 6103
rect 13084 6060 13136 6069
rect 15476 6060 15528 6112
rect 16488 6103 16540 6112
rect 16488 6069 16497 6103
rect 16497 6069 16531 6103
rect 16531 6069 16540 6103
rect 16488 6060 16540 6069
rect 16856 6060 16908 6112
rect 18052 6060 18104 6112
rect 19340 6060 19392 6112
rect 20628 6060 20680 6112
rect 21180 6060 21232 6112
rect 3595 5958 3647 6010
rect 3659 5958 3711 6010
rect 3723 5958 3775 6010
rect 3787 5958 3839 6010
rect 3851 5958 3903 6010
rect 8885 5958 8937 6010
rect 8949 5958 9001 6010
rect 9013 5958 9065 6010
rect 9077 5958 9129 6010
rect 9141 5958 9193 6010
rect 14175 5958 14227 6010
rect 14239 5958 14291 6010
rect 14303 5958 14355 6010
rect 14367 5958 14419 6010
rect 14431 5958 14483 6010
rect 19465 5958 19517 6010
rect 19529 5958 19581 6010
rect 19593 5958 19645 6010
rect 19657 5958 19709 6010
rect 19721 5958 19773 6010
rect 3240 5856 3292 5908
rect 3976 5652 4028 5704
rect 4160 5652 4212 5704
rect 4620 5584 4672 5636
rect 6276 5831 6328 5840
rect 6276 5797 6285 5831
rect 6285 5797 6319 5831
rect 6319 5797 6328 5831
rect 6276 5788 6328 5797
rect 7564 5856 7616 5908
rect 7288 5788 7340 5840
rect 5540 5720 5592 5772
rect 8576 5856 8628 5908
rect 9404 5856 9456 5908
rect 9772 5899 9824 5908
rect 9772 5865 9781 5899
rect 9781 5865 9815 5899
rect 9815 5865 9824 5899
rect 9772 5856 9824 5865
rect 9956 5856 10008 5908
rect 13084 5856 13136 5908
rect 15476 5899 15528 5908
rect 15476 5865 15485 5899
rect 15485 5865 15519 5899
rect 15519 5865 15528 5899
rect 15476 5856 15528 5865
rect 16028 5899 16080 5908
rect 16028 5865 16037 5899
rect 16037 5865 16071 5899
rect 16071 5865 16080 5899
rect 16028 5856 16080 5865
rect 16488 5856 16540 5908
rect 20260 5899 20312 5908
rect 20260 5865 20269 5899
rect 20269 5865 20303 5899
rect 20303 5865 20312 5899
rect 20260 5856 20312 5865
rect 6460 5627 6512 5636
rect 5632 5516 5684 5568
rect 6460 5593 6487 5627
rect 6487 5593 6512 5627
rect 6460 5584 6512 5593
rect 6920 5652 6972 5704
rect 9220 5720 9272 5772
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 8668 5652 8720 5704
rect 8024 5627 8076 5636
rect 8024 5593 8064 5627
rect 8064 5593 8076 5627
rect 8024 5584 8076 5593
rect 8668 5516 8720 5568
rect 8852 5652 8904 5704
rect 9220 5584 9272 5636
rect 9312 5584 9364 5636
rect 9680 5584 9732 5636
rect 9404 5516 9456 5568
rect 9864 5695 9916 5704
rect 9864 5661 9873 5695
rect 9873 5661 9907 5695
rect 9907 5661 9916 5695
rect 9864 5652 9916 5661
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 10600 5763 10652 5772
rect 10600 5729 10609 5763
rect 10609 5729 10643 5763
rect 10643 5729 10652 5763
rect 10600 5720 10652 5729
rect 11152 5695 11204 5704
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 11152 5652 11204 5661
rect 12072 5652 12124 5704
rect 19892 5720 19944 5772
rect 21180 5763 21232 5772
rect 21180 5729 21189 5763
rect 21189 5729 21223 5763
rect 21223 5729 21232 5763
rect 21180 5720 21232 5729
rect 13268 5652 13320 5704
rect 13728 5652 13780 5704
rect 15292 5652 15344 5704
rect 16856 5652 16908 5704
rect 18144 5652 18196 5704
rect 20536 5652 20588 5704
rect 12164 5627 12216 5636
rect 12164 5593 12173 5627
rect 12173 5593 12207 5627
rect 12207 5593 12216 5627
rect 12164 5584 12216 5593
rect 13820 5584 13872 5636
rect 18052 5559 18104 5568
rect 18052 5525 18061 5559
rect 18061 5525 18095 5559
rect 18095 5525 18104 5559
rect 18052 5516 18104 5525
rect 19892 5516 19944 5568
rect 20628 5559 20680 5568
rect 20628 5525 20637 5559
rect 20637 5525 20671 5559
rect 20671 5525 20680 5559
rect 20628 5516 20680 5525
rect 4255 5414 4307 5466
rect 4319 5414 4371 5466
rect 4383 5414 4435 5466
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 9545 5414 9597 5466
rect 9609 5414 9661 5466
rect 9673 5414 9725 5466
rect 9737 5414 9789 5466
rect 9801 5414 9853 5466
rect 14835 5414 14887 5466
rect 14899 5414 14951 5466
rect 14963 5414 15015 5466
rect 15027 5414 15079 5466
rect 15091 5414 15143 5466
rect 20125 5414 20177 5466
rect 20189 5414 20241 5466
rect 20253 5414 20305 5466
rect 20317 5414 20369 5466
rect 20381 5414 20433 5466
rect 4620 5312 4672 5364
rect 7564 5312 7616 5364
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 5080 5219 5132 5228
rect 5080 5185 5089 5219
rect 5089 5185 5123 5219
rect 5123 5185 5132 5219
rect 5080 5176 5132 5185
rect 6920 5244 6972 5296
rect 5632 5176 5684 5228
rect 5816 5176 5868 5228
rect 6092 5176 6144 5228
rect 7104 5176 7156 5228
rect 7472 5176 7524 5228
rect 10600 5312 10652 5364
rect 14648 5312 14700 5364
rect 19340 5312 19392 5364
rect 19984 5312 20036 5364
rect 20536 5312 20588 5364
rect 20720 5312 20772 5364
rect 21824 5312 21876 5364
rect 14740 5287 14792 5296
rect 14740 5253 14749 5287
rect 14749 5253 14783 5287
rect 14783 5253 14792 5287
rect 14740 5244 14792 5253
rect 9312 5176 9364 5228
rect 9864 5176 9916 5228
rect 10048 5176 10100 5228
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 16396 5176 16448 5228
rect 17132 5176 17184 5228
rect 18052 5176 18104 5228
rect 19892 5176 19944 5228
rect 20628 5219 20680 5228
rect 20628 5185 20637 5219
rect 20637 5185 20671 5219
rect 20671 5185 20680 5219
rect 20628 5176 20680 5185
rect 7748 5108 7800 5160
rect 16304 5151 16356 5160
rect 16304 5117 16313 5151
rect 16313 5117 16347 5151
rect 16347 5117 16356 5151
rect 16304 5108 16356 5117
rect 1860 4972 1912 5024
rect 7564 5015 7616 5024
rect 7564 4981 7573 5015
rect 7573 4981 7607 5015
rect 7607 4981 7616 5015
rect 7564 4972 7616 4981
rect 7656 4972 7708 5024
rect 12900 4972 12952 5024
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 15384 4972 15436 5024
rect 17224 4972 17276 5024
rect 3595 4870 3647 4922
rect 3659 4870 3711 4922
rect 3723 4870 3775 4922
rect 3787 4870 3839 4922
rect 3851 4870 3903 4922
rect 8885 4870 8937 4922
rect 8949 4870 9001 4922
rect 9013 4870 9065 4922
rect 9077 4870 9129 4922
rect 9141 4870 9193 4922
rect 14175 4870 14227 4922
rect 14239 4870 14291 4922
rect 14303 4870 14355 4922
rect 14367 4870 14419 4922
rect 14431 4870 14483 4922
rect 19465 4870 19517 4922
rect 19529 4870 19581 4922
rect 19593 4870 19645 4922
rect 19657 4870 19709 4922
rect 19721 4870 19773 4922
rect 4804 4564 4856 4616
rect 5080 4564 5132 4616
rect 6276 4768 6328 4820
rect 7564 4768 7616 4820
rect 7656 4768 7708 4820
rect 13728 4768 13780 4820
rect 13820 4811 13872 4820
rect 13820 4777 13829 4811
rect 13829 4777 13863 4811
rect 13863 4777 13872 4811
rect 13820 4768 13872 4777
rect 15752 4768 15804 4820
rect 16028 4768 16080 4820
rect 16304 4768 16356 4820
rect 7472 4700 7524 4752
rect 5908 4632 5960 4684
rect 7748 4700 7800 4752
rect 11704 4700 11756 4752
rect 7656 4675 7708 4684
rect 7656 4641 7665 4675
rect 7665 4641 7699 4675
rect 7699 4641 7708 4675
rect 7656 4632 7708 4641
rect 5356 4539 5408 4548
rect 5356 4505 5365 4539
rect 5365 4505 5399 4539
rect 5399 4505 5408 4539
rect 6092 4564 6144 4616
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 7380 4564 7432 4616
rect 15200 4632 15252 4684
rect 13636 4607 13688 4616
rect 13636 4573 13645 4607
rect 13645 4573 13679 4607
rect 13679 4573 13688 4607
rect 13636 4564 13688 4573
rect 15384 4564 15436 4616
rect 15660 4607 15712 4616
rect 15660 4573 15669 4607
rect 15669 4573 15703 4607
rect 15703 4573 15712 4607
rect 15660 4564 15712 4573
rect 16672 4564 16724 4616
rect 17224 4768 17276 4820
rect 17868 4564 17920 4616
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 5356 4496 5408 4505
rect 16856 4496 16908 4548
rect 5632 4428 5684 4480
rect 8116 4428 8168 4480
rect 13728 4428 13780 4480
rect 16212 4428 16264 4480
rect 18420 4471 18472 4480
rect 18420 4437 18429 4471
rect 18429 4437 18463 4471
rect 18463 4437 18472 4471
rect 18420 4428 18472 4437
rect 18696 4471 18748 4480
rect 18696 4437 18705 4471
rect 18705 4437 18739 4471
rect 18739 4437 18748 4471
rect 18696 4428 18748 4437
rect 4255 4326 4307 4378
rect 4319 4326 4371 4378
rect 4383 4326 4435 4378
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 9545 4326 9597 4378
rect 9609 4326 9661 4378
rect 9673 4326 9725 4378
rect 9737 4326 9789 4378
rect 9801 4326 9853 4378
rect 14835 4326 14887 4378
rect 14899 4326 14951 4378
rect 14963 4326 15015 4378
rect 15027 4326 15079 4378
rect 15091 4326 15143 4378
rect 20125 4326 20177 4378
rect 20189 4326 20241 4378
rect 20253 4326 20305 4378
rect 20317 4326 20369 4378
rect 20381 4326 20433 4378
rect 7932 4156 7984 4208
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 5632 4020 5684 4072
rect 5908 4020 5960 4072
rect 8024 4088 8076 4140
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 4620 3884 4672 3936
rect 5080 3884 5132 3936
rect 6828 3884 6880 3936
rect 6920 3884 6972 3936
rect 8208 3884 8260 3936
rect 8484 3884 8536 3936
rect 8668 4088 8720 4140
rect 9772 4156 9824 4208
rect 11704 4224 11756 4276
rect 15200 4267 15252 4276
rect 15200 4233 15209 4267
rect 15209 4233 15243 4267
rect 15243 4233 15252 4267
rect 15200 4224 15252 4233
rect 15384 4224 15436 4276
rect 16672 4267 16724 4276
rect 16672 4233 16681 4267
rect 16681 4233 16715 4267
rect 16715 4233 16724 4267
rect 16672 4224 16724 4233
rect 17684 4224 17736 4276
rect 17868 4224 17920 4276
rect 18420 4224 18472 4276
rect 19984 4224 20036 4276
rect 12624 4156 12676 4208
rect 13728 4156 13780 4208
rect 9220 4088 9272 4140
rect 9588 4131 9640 4140
rect 9588 4097 9597 4131
rect 9597 4097 9631 4131
rect 9631 4097 9640 4131
rect 9588 4088 9640 4097
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 11704 4088 11756 4140
rect 16120 4199 16172 4208
rect 16120 4165 16145 4199
rect 16145 4165 16172 4199
rect 16120 4156 16172 4165
rect 16488 4156 16540 4208
rect 9588 3952 9640 4004
rect 10692 3884 10744 3936
rect 11060 3884 11112 3936
rect 11704 3995 11756 4004
rect 11704 3961 11713 3995
rect 11713 3961 11747 3995
rect 11747 3961 11756 3995
rect 11704 3952 11756 3961
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 12900 3884 12952 3936
rect 17040 4199 17092 4208
rect 17040 4165 17049 4199
rect 17049 4165 17083 4199
rect 17083 4165 17092 4199
rect 17040 4156 17092 4165
rect 18696 4156 18748 4208
rect 13452 3927 13504 3936
rect 13452 3893 13461 3927
rect 13461 3893 13495 3927
rect 13495 3893 13504 3927
rect 13452 3884 13504 3893
rect 14740 3884 14792 3936
rect 16580 3884 16632 3936
rect 19340 4088 19392 4140
rect 20168 4088 20220 4140
rect 18052 4020 18104 4072
rect 17776 3884 17828 3936
rect 18144 3884 18196 3936
rect 19800 3884 19852 3936
rect 3595 3782 3647 3834
rect 3659 3782 3711 3834
rect 3723 3782 3775 3834
rect 3787 3782 3839 3834
rect 3851 3782 3903 3834
rect 8885 3782 8937 3834
rect 8949 3782 9001 3834
rect 9013 3782 9065 3834
rect 9077 3782 9129 3834
rect 9141 3782 9193 3834
rect 14175 3782 14227 3834
rect 14239 3782 14291 3834
rect 14303 3782 14355 3834
rect 14367 3782 14419 3834
rect 14431 3782 14483 3834
rect 19465 3782 19517 3834
rect 19529 3782 19581 3834
rect 19593 3782 19645 3834
rect 19657 3782 19709 3834
rect 19721 3782 19773 3834
rect 7288 3680 7340 3732
rect 6920 3612 6972 3664
rect 8392 3680 8444 3732
rect 8024 3612 8076 3664
rect 9588 3612 9640 3664
rect 5540 3476 5592 3528
rect 7932 3476 7984 3528
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 5080 3408 5132 3460
rect 6828 3408 6880 3460
rect 8668 3544 8720 3596
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 9220 3476 9272 3528
rect 9772 3680 9824 3732
rect 11244 3680 11296 3732
rect 10692 3655 10744 3664
rect 10692 3621 10701 3655
rect 10701 3621 10735 3655
rect 10735 3621 10744 3655
rect 10692 3612 10744 3621
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12440 3680 12492 3689
rect 12624 3680 12676 3732
rect 13636 3680 13688 3732
rect 15660 3680 15712 3732
rect 16488 3723 16540 3732
rect 16488 3689 16497 3723
rect 16497 3689 16531 3723
rect 16531 3689 16540 3723
rect 16488 3680 16540 3689
rect 16856 3680 16908 3732
rect 17868 3723 17920 3732
rect 17868 3689 17877 3723
rect 17877 3689 17911 3723
rect 17911 3689 17920 3723
rect 17868 3680 17920 3689
rect 10508 3476 10560 3528
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 10876 3476 10928 3528
rect 11152 3476 11204 3528
rect 8484 3340 8536 3392
rect 9404 3340 9456 3392
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 12072 3476 12124 3485
rect 12164 3476 12216 3528
rect 17960 3612 18012 3664
rect 12900 3544 12952 3596
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 16396 3544 16448 3596
rect 12992 3519 13044 3528
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 12992 3476 13044 3485
rect 13176 3519 13228 3528
rect 13176 3485 13185 3519
rect 13185 3485 13219 3519
rect 13219 3485 13228 3519
rect 13176 3476 13228 3485
rect 13452 3476 13504 3528
rect 13728 3476 13780 3528
rect 10048 3383 10100 3392
rect 10048 3349 10057 3383
rect 10057 3349 10091 3383
rect 10091 3349 10100 3383
rect 10048 3340 10100 3349
rect 10416 3340 10468 3392
rect 10876 3383 10928 3392
rect 10876 3349 10885 3383
rect 10885 3349 10919 3383
rect 10919 3349 10928 3383
rect 16580 3519 16632 3528
rect 16580 3485 16589 3519
rect 16589 3485 16623 3519
rect 16623 3485 16632 3519
rect 16580 3476 16632 3485
rect 18512 3680 18564 3732
rect 20168 3723 20220 3732
rect 20168 3689 20177 3723
rect 20177 3689 20211 3723
rect 20211 3689 20220 3723
rect 20168 3680 20220 3689
rect 17040 3476 17092 3528
rect 17132 3519 17184 3528
rect 17132 3485 17141 3519
rect 17141 3485 17175 3519
rect 17175 3485 17184 3519
rect 17132 3476 17184 3485
rect 16672 3408 16724 3460
rect 17776 3476 17828 3528
rect 18144 3476 18196 3528
rect 19800 3519 19852 3528
rect 19800 3485 19809 3519
rect 19809 3485 19843 3519
rect 19843 3485 19852 3519
rect 19800 3476 19852 3485
rect 19984 3519 20036 3528
rect 19984 3485 19993 3519
rect 19993 3485 20027 3519
rect 20027 3485 20036 3519
rect 19984 3476 20036 3485
rect 10876 3340 10928 3349
rect 13268 3340 13320 3392
rect 13452 3383 13504 3392
rect 13452 3349 13461 3383
rect 13461 3349 13495 3383
rect 13495 3349 13504 3383
rect 13452 3340 13504 3349
rect 17868 3451 17920 3460
rect 17868 3417 17877 3451
rect 17877 3417 17911 3451
rect 17911 3417 17920 3451
rect 17868 3408 17920 3417
rect 18052 3340 18104 3392
rect 18512 3340 18564 3392
rect 4255 3238 4307 3290
rect 4319 3238 4371 3290
rect 4383 3238 4435 3290
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 9545 3238 9597 3290
rect 9609 3238 9661 3290
rect 9673 3238 9725 3290
rect 9737 3238 9789 3290
rect 9801 3238 9853 3290
rect 14835 3238 14887 3290
rect 14899 3238 14951 3290
rect 14963 3238 15015 3290
rect 15027 3238 15079 3290
rect 15091 3238 15143 3290
rect 20125 3238 20177 3290
rect 20189 3238 20241 3290
rect 20253 3238 20305 3290
rect 20317 3238 20369 3290
rect 20381 3238 20433 3290
rect 4620 3136 4672 3188
rect 5172 3136 5224 3188
rect 6092 3136 6144 3188
rect 6276 3136 6328 3188
rect 6828 3179 6880 3188
rect 4160 3000 4212 3052
rect 6828 3145 6837 3179
rect 6837 3145 6871 3179
rect 6871 3145 6880 3179
rect 6828 3136 6880 3145
rect 6920 3136 6972 3188
rect 8208 3136 8260 3188
rect 8300 3136 8352 3188
rect 5908 2864 5960 2916
rect 6276 2864 6328 2916
rect 8484 3000 8536 3052
rect 10048 3136 10100 3188
rect 11152 3136 11204 3188
rect 10784 3068 10836 3120
rect 9496 3000 9548 3052
rect 11060 3043 11112 3052
rect 11060 3009 11081 3043
rect 11081 3009 11112 3043
rect 11060 3000 11112 3009
rect 11244 3000 11296 3052
rect 12440 3136 12492 3188
rect 14740 3136 14792 3188
rect 11796 3068 11848 3120
rect 12072 3068 12124 3120
rect 11612 3000 11664 3052
rect 6552 2839 6604 2848
rect 6552 2805 6561 2839
rect 6561 2805 6595 2839
rect 6595 2805 6604 2839
rect 6552 2796 6604 2805
rect 10600 2864 10652 2916
rect 10876 2864 10928 2916
rect 12900 3043 12952 3052
rect 12900 3009 12909 3043
rect 12909 3009 12943 3043
rect 12943 3009 12952 3043
rect 12900 3000 12952 3009
rect 13176 3043 13228 3052
rect 13176 3009 13210 3043
rect 13210 3009 13228 3043
rect 13176 3000 13228 3009
rect 16212 3136 16264 3188
rect 16396 3136 16448 3188
rect 17132 3136 17184 3188
rect 18144 3136 18196 3188
rect 19340 3136 19392 3188
rect 19984 3136 20036 3188
rect 17500 3000 17552 3052
rect 18880 3000 18932 3052
rect 21456 3000 21508 3052
rect 16672 2932 16724 2984
rect 12164 2907 12216 2916
rect 12164 2873 12173 2907
rect 12173 2873 12207 2907
rect 12207 2873 12216 2907
rect 12164 2864 12216 2873
rect 8024 2796 8076 2848
rect 8576 2839 8628 2848
rect 8576 2805 8585 2839
rect 8585 2805 8619 2839
rect 8619 2805 8628 2839
rect 8576 2796 8628 2805
rect 9220 2796 9272 2848
rect 11612 2796 11664 2848
rect 13268 2796 13320 2848
rect 18512 2796 18564 2848
rect 3595 2694 3647 2746
rect 3659 2694 3711 2746
rect 3723 2694 3775 2746
rect 3787 2694 3839 2746
rect 3851 2694 3903 2746
rect 8885 2694 8937 2746
rect 8949 2694 9001 2746
rect 9013 2694 9065 2746
rect 9077 2694 9129 2746
rect 9141 2694 9193 2746
rect 14175 2694 14227 2746
rect 14239 2694 14291 2746
rect 14303 2694 14355 2746
rect 14367 2694 14419 2746
rect 14431 2694 14483 2746
rect 19465 2694 19517 2746
rect 19529 2694 19581 2746
rect 19593 2694 19645 2746
rect 19657 2694 19709 2746
rect 19721 2694 19773 2746
rect 13176 2592 13228 2644
rect 17500 2592 17552 2644
rect 17960 2592 18012 2644
rect 18880 2635 18932 2644
rect 18880 2601 18889 2635
rect 18889 2601 18923 2635
rect 18923 2601 18932 2635
rect 18880 2592 18932 2601
rect 18972 2592 19024 2644
rect 21456 2635 21508 2644
rect 21456 2601 21465 2635
rect 21465 2601 21499 2635
rect 21499 2601 21508 2635
rect 21456 2592 21508 2601
rect 17132 2456 17184 2508
rect 20 2388 72 2440
rect 8576 2388 8628 2440
rect 13544 2431 13596 2440
rect 13544 2397 13553 2431
rect 13553 2397 13587 2431
rect 13587 2397 13596 2431
rect 13544 2388 13596 2397
rect 18512 2499 18564 2508
rect 18512 2465 18521 2499
rect 18521 2465 18555 2499
rect 18555 2465 18564 2499
rect 18512 2456 18564 2465
rect 17868 2320 17920 2372
rect 8392 2252 8444 2304
rect 13084 2252 13136 2304
rect 22192 2252 22244 2304
rect 4255 2150 4307 2202
rect 4319 2150 4371 2202
rect 4383 2150 4435 2202
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 9545 2150 9597 2202
rect 9609 2150 9661 2202
rect 9673 2150 9725 2202
rect 9737 2150 9789 2202
rect 9801 2150 9853 2202
rect 14835 2150 14887 2202
rect 14899 2150 14951 2202
rect 14963 2150 15015 2202
rect 15027 2150 15079 2202
rect 15091 2150 15143 2202
rect 20125 2150 20177 2202
rect 20189 2150 20241 2202
rect 20253 2150 20305 2202
rect 20317 2150 20369 2202
rect 20381 2150 20433 2202
<< metal2 >>
rect 1306 24752 1362 25552
rect 10322 24752 10378 25552
rect 19338 24752 19394 25552
rect 1320 22778 1348 24752
rect 4255 22876 4563 22885
rect 4255 22874 4261 22876
rect 4317 22874 4341 22876
rect 4397 22874 4421 22876
rect 4477 22874 4501 22876
rect 4557 22874 4563 22876
rect 4317 22822 4319 22874
rect 4499 22822 4501 22874
rect 4255 22820 4261 22822
rect 4317 22820 4341 22822
rect 4397 22820 4421 22822
rect 4477 22820 4501 22822
rect 4557 22820 4563 22822
rect 4255 22811 4563 22820
rect 9545 22876 9853 22885
rect 9545 22874 9551 22876
rect 9607 22874 9631 22876
rect 9687 22874 9711 22876
rect 9767 22874 9791 22876
rect 9847 22874 9853 22876
rect 9607 22822 9609 22874
rect 9789 22822 9791 22874
rect 9545 22820 9551 22822
rect 9607 22820 9631 22822
rect 9687 22820 9711 22822
rect 9767 22820 9791 22822
rect 9847 22820 9853 22822
rect 9545 22811 9853 22820
rect 10336 22778 10364 24752
rect 14835 22876 15143 22885
rect 14835 22874 14841 22876
rect 14897 22874 14921 22876
rect 14977 22874 15001 22876
rect 15057 22874 15081 22876
rect 15137 22874 15143 22876
rect 14897 22822 14899 22874
rect 15079 22822 15081 22874
rect 14835 22820 14841 22822
rect 14897 22820 14921 22822
rect 14977 22820 15001 22822
rect 15057 22820 15081 22822
rect 15137 22820 15143 22822
rect 14835 22811 15143 22820
rect 19352 22778 19380 24752
rect 20125 22876 20433 22885
rect 20125 22874 20131 22876
rect 20187 22874 20211 22876
rect 20267 22874 20291 22876
rect 20347 22874 20371 22876
rect 20427 22874 20433 22876
rect 20187 22822 20189 22874
rect 20369 22822 20371 22874
rect 20125 22820 20131 22822
rect 20187 22820 20211 22822
rect 20267 22820 20291 22822
rect 20347 22820 20371 22822
rect 20427 22820 20433 22822
rect 20125 22811 20433 22820
rect 1308 22772 1360 22778
rect 1308 22714 1360 22720
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 1780 21486 1808 22578
rect 3595 22332 3903 22341
rect 3595 22330 3601 22332
rect 3657 22330 3681 22332
rect 3737 22330 3761 22332
rect 3817 22330 3841 22332
rect 3897 22330 3903 22332
rect 3657 22278 3659 22330
rect 3839 22278 3841 22330
rect 3595 22276 3601 22278
rect 3657 22276 3681 22278
rect 3737 22276 3761 22278
rect 3817 22276 3841 22278
rect 3897 22276 3903 22278
rect 3595 22267 3903 22276
rect 8885 22332 9193 22341
rect 8885 22330 8891 22332
rect 8947 22330 8971 22332
rect 9027 22330 9051 22332
rect 9107 22330 9131 22332
rect 9187 22330 9193 22332
rect 8947 22278 8949 22330
rect 9129 22278 9131 22330
rect 8885 22276 8891 22278
rect 8947 22276 8971 22278
rect 9027 22276 9051 22278
rect 9107 22276 9131 22278
rect 9187 22276 9193 22278
rect 8885 22267 9193 22276
rect 7564 22160 7616 22166
rect 7564 22102 7616 22108
rect 8392 22160 8444 22166
rect 8392 22102 8444 22108
rect 12992 22160 13044 22166
rect 12992 22102 13044 22108
rect 2596 22092 2648 22098
rect 2596 22034 2648 22040
rect 4896 22092 4948 22098
rect 4896 22034 4948 22040
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 1768 21480 1820 21486
rect 1768 21422 1820 21428
rect 2516 21146 2544 21490
rect 2608 21418 2636 22034
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 2964 21956 3016 21962
rect 2964 21898 3016 21904
rect 2596 21412 2648 21418
rect 2596 21354 2648 21360
rect 2504 21140 2556 21146
rect 2504 21082 2556 21088
rect 2608 19446 2636 21354
rect 2976 21146 3004 21898
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 3068 21690 3096 21830
rect 3056 21684 3108 21690
rect 3056 21626 3108 21632
rect 3436 21146 3464 21966
rect 3516 21888 3568 21894
rect 3516 21830 3568 21836
rect 4068 21888 4120 21894
rect 4068 21830 4120 21836
rect 3528 21146 3556 21830
rect 4080 21418 4108 21830
rect 4255 21788 4563 21797
rect 4255 21786 4261 21788
rect 4317 21786 4341 21788
rect 4397 21786 4421 21788
rect 4477 21786 4501 21788
rect 4557 21786 4563 21788
rect 4317 21734 4319 21786
rect 4499 21734 4501 21786
rect 4255 21732 4261 21734
rect 4317 21732 4341 21734
rect 4397 21732 4421 21734
rect 4477 21732 4501 21734
rect 4557 21732 4563 21734
rect 4255 21723 4563 21732
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 3595 21244 3903 21253
rect 3595 21242 3601 21244
rect 3657 21242 3681 21244
rect 3737 21242 3761 21244
rect 3817 21242 3841 21244
rect 3897 21242 3903 21244
rect 3657 21190 3659 21242
rect 3839 21190 3841 21242
rect 3595 21188 3601 21190
rect 3657 21188 3681 21190
rect 3737 21188 3761 21190
rect 3817 21188 3841 21190
rect 3897 21188 3903 21190
rect 3595 21179 3903 21188
rect 3988 21146 4016 21286
rect 4080 21146 4108 21354
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 3148 20936 3200 20942
rect 3148 20878 3200 20884
rect 3160 20262 3188 20878
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 2596 19440 2648 19446
rect 2596 19382 2648 19388
rect 2608 18970 2636 19382
rect 2596 18964 2648 18970
rect 2596 18906 2648 18912
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2792 18426 2820 18634
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2976 18290 3004 19654
rect 3068 19378 3096 19654
rect 3056 19372 3108 19378
rect 3056 19314 3108 19320
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1504 16658 1532 17138
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1504 15026 1532 16594
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1688 16250 1716 16390
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 2148 16182 2176 16458
rect 2136 16176 2188 16182
rect 2136 16118 2188 16124
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2332 15706 2360 16050
rect 2320 15700 2372 15706
rect 3160 15688 3188 20198
rect 3436 19854 3464 21082
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3988 20602 4016 20878
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3976 20324 4028 20330
rect 3976 20266 4028 20272
rect 3595 20156 3903 20165
rect 3595 20154 3601 20156
rect 3657 20154 3681 20156
rect 3737 20154 3761 20156
rect 3817 20154 3841 20156
rect 3897 20154 3903 20156
rect 3657 20102 3659 20154
rect 3839 20102 3841 20154
rect 3595 20100 3601 20102
rect 3657 20100 3681 20102
rect 3737 20100 3761 20102
rect 3817 20100 3841 20102
rect 3897 20100 3903 20102
rect 3595 20091 3903 20100
rect 3988 19854 4016 20266
rect 3240 19848 3292 19854
rect 3424 19848 3476 19854
rect 3240 19790 3292 19796
rect 3344 19796 3424 19802
rect 3344 19790 3476 19796
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3252 19378 3280 19790
rect 3344 19774 3464 19790
rect 3344 19514 3372 19774
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3436 19378 3464 19654
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3344 18086 3372 19110
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3344 17678 3372 18022
rect 3528 17678 3556 19790
rect 3988 19514 4016 19790
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3595 19068 3903 19077
rect 3595 19066 3601 19068
rect 3657 19066 3681 19068
rect 3737 19066 3761 19068
rect 3817 19066 3841 19068
rect 3897 19066 3903 19068
rect 3657 19014 3659 19066
rect 3839 19014 3841 19066
rect 3595 19012 3601 19014
rect 3657 19012 3681 19014
rect 3737 19012 3761 19014
rect 3817 19012 3841 19014
rect 3897 19012 3903 19014
rect 3595 19003 3903 19012
rect 3988 18630 4016 19110
rect 4080 18970 4108 20878
rect 4255 20700 4563 20709
rect 4255 20698 4261 20700
rect 4317 20698 4341 20700
rect 4397 20698 4421 20700
rect 4477 20698 4501 20700
rect 4557 20698 4563 20700
rect 4317 20646 4319 20698
rect 4499 20646 4501 20698
rect 4255 20644 4261 20646
rect 4317 20644 4341 20646
rect 4397 20644 4421 20646
rect 4477 20644 4501 20646
rect 4557 20644 4563 20646
rect 4255 20635 4563 20644
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4255 19612 4563 19621
rect 4255 19610 4261 19612
rect 4317 19610 4341 19612
rect 4397 19610 4421 19612
rect 4477 19610 4501 19612
rect 4557 19610 4563 19612
rect 4317 19558 4319 19610
rect 4499 19558 4501 19610
rect 4255 19556 4261 19558
rect 4317 19556 4341 19558
rect 4397 19556 4421 19558
rect 4477 19556 4501 19558
rect 4557 19556 4563 19558
rect 4255 19547 4563 19556
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4632 18766 4660 19654
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4620 18624 4672 18630
rect 4620 18566 4672 18572
rect 3988 18222 4016 18566
rect 4172 18426 4200 18566
rect 4255 18524 4563 18533
rect 4255 18522 4261 18524
rect 4317 18522 4341 18524
rect 4397 18522 4421 18524
rect 4477 18522 4501 18524
rect 4557 18522 4563 18524
rect 4317 18470 4319 18522
rect 4499 18470 4501 18522
rect 4255 18468 4261 18470
rect 4317 18468 4341 18470
rect 4397 18468 4421 18470
rect 4477 18468 4501 18470
rect 4557 18468 4563 18470
rect 4255 18459 4563 18468
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4528 18284 4580 18290
rect 4528 18226 4580 18232
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3595 17980 3903 17989
rect 3595 17978 3601 17980
rect 3657 17978 3681 17980
rect 3737 17978 3761 17980
rect 3817 17978 3841 17980
rect 3897 17978 3903 17980
rect 3657 17926 3659 17978
rect 3839 17926 3841 17978
rect 3595 17924 3601 17926
rect 3657 17924 3681 17926
rect 3737 17924 3761 17926
rect 3817 17924 3841 17926
rect 3897 17924 3903 17926
rect 3595 17915 3903 17924
rect 4540 17746 4568 18226
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4528 17740 4580 17746
rect 4528 17682 4580 17688
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3252 16114 3280 16934
rect 3344 16726 3372 17614
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3528 17338 3556 17478
rect 3804 17338 3832 17478
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3608 17196 3660 17202
rect 3528 17156 3608 17184
rect 3332 16720 3384 16726
rect 3332 16662 3384 16668
rect 3528 16590 3556 17156
rect 3608 17138 3660 17144
rect 4080 17066 4108 17682
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4172 17202 4200 17478
rect 4255 17436 4563 17445
rect 4255 17434 4261 17436
rect 4317 17434 4341 17436
rect 4397 17434 4421 17436
rect 4477 17434 4501 17436
rect 4557 17434 4563 17436
rect 4317 17382 4319 17434
rect 4499 17382 4501 17434
rect 4255 17380 4261 17382
rect 4317 17380 4341 17382
rect 4397 17380 4421 17382
rect 4477 17380 4501 17382
rect 4557 17380 4563 17382
rect 4255 17371 4563 17380
rect 4632 17338 4660 18566
rect 4724 18426 4752 18770
rect 4816 18426 4844 19654
rect 4908 18834 4936 22034
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 5724 21956 5776 21962
rect 5724 21898 5776 21904
rect 5736 21690 5764 21898
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 6092 21616 6144 21622
rect 6092 21558 6144 21564
rect 5724 21412 5776 21418
rect 5776 21372 5856 21400
rect 5724 21354 5776 21360
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5552 21010 5580 21286
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5828 20942 5856 21372
rect 6104 21010 6132 21558
rect 6748 21554 6776 21966
rect 7380 21956 7432 21962
rect 7380 21898 7432 21904
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6196 21146 6224 21490
rect 6276 21480 6328 21486
rect 6748 21457 6776 21490
rect 6276 21422 6328 21428
rect 6734 21448 6790 21457
rect 6288 21146 6316 21422
rect 6734 21383 6790 21392
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6736 21344 6788 21350
rect 6736 21286 6788 21292
rect 6184 21140 6236 21146
rect 6184 21082 6236 21088
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6656 21010 6684 21286
rect 6748 21146 6776 21286
rect 6840 21146 6868 21626
rect 7116 21554 7144 21830
rect 7208 21690 7236 21830
rect 7196 21684 7248 21690
rect 7196 21626 7248 21632
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 5828 20806 5856 20878
rect 5816 20800 5868 20806
rect 5816 20742 5868 20748
rect 5920 20602 5948 20878
rect 6656 20618 6684 20946
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 5908 20596 5960 20602
rect 6656 20590 6776 20618
rect 5908 20538 5960 20544
rect 6748 20466 6776 20590
rect 6840 20466 6868 20742
rect 6932 20602 6960 21422
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 7116 20602 7144 21286
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 7104 20596 7156 20602
rect 7208 20584 7236 21626
rect 7392 21146 7420 21898
rect 7576 21486 7604 22102
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7654 21448 7710 21457
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7576 20942 7604 21422
rect 7654 21383 7710 21392
rect 7668 20942 7696 21383
rect 7760 21146 7788 21830
rect 7852 21622 7880 21830
rect 7840 21616 7892 21622
rect 7840 21558 7892 21564
rect 7852 21146 7880 21558
rect 8312 21146 8340 21966
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 8300 21140 8352 21146
rect 8404 21128 8432 22102
rect 12716 22092 12768 22098
rect 12716 22034 12768 22040
rect 9956 22024 10008 22030
rect 12072 22024 12124 22030
rect 9956 21966 10008 21972
rect 11992 21972 12072 21978
rect 11992 21966 12124 21972
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8496 21622 8524 21830
rect 9545 21788 9853 21797
rect 9545 21786 9551 21788
rect 9607 21786 9631 21788
rect 9687 21786 9711 21788
rect 9767 21786 9791 21788
rect 9847 21786 9853 21788
rect 9607 21734 9609 21786
rect 9789 21734 9791 21786
rect 9545 21732 9551 21734
rect 9607 21732 9631 21734
rect 9687 21732 9711 21734
rect 9767 21732 9791 21734
rect 9847 21732 9853 21734
rect 9545 21723 9853 21732
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 9864 21344 9916 21350
rect 9968 21332 9996 21966
rect 10416 21956 10468 21962
rect 10416 21898 10468 21904
rect 11992 21950 12112 21966
rect 12164 21956 12216 21962
rect 10428 21690 10456 21898
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 11440 21690 11468 21830
rect 11992 21706 12020 21950
rect 12164 21898 12216 21904
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 11900 21690 12020 21706
rect 12084 21690 12112 21830
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 11888 21684 12020 21690
rect 11940 21678 12020 21684
rect 11888 21626 11940 21632
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 9916 21304 9996 21332
rect 10784 21344 10836 21350
rect 9864 21286 9916 21292
rect 10784 21286 10836 21292
rect 8885 21244 9193 21253
rect 8885 21242 8891 21244
rect 8947 21242 8971 21244
rect 9027 21242 9051 21244
rect 9107 21242 9131 21244
rect 9187 21242 9193 21244
rect 8947 21190 8949 21242
rect 9129 21190 9131 21242
rect 8885 21188 8891 21190
rect 8947 21188 8971 21190
rect 9027 21188 9051 21190
rect 9107 21188 9131 21190
rect 9187 21188 9193 21190
rect 8885 21179 9193 21188
rect 8484 21140 8536 21146
rect 8404 21100 8484 21128
rect 8300 21082 8352 21088
rect 8484 21082 8536 21088
rect 9876 20942 9904 21286
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 9864 20936 9916 20942
rect 9916 20896 9996 20924
rect 9864 20878 9916 20884
rect 7288 20596 7340 20602
rect 7208 20556 7288 20584
rect 7104 20538 7156 20544
rect 7288 20538 7340 20544
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6748 19854 6776 20402
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6840 19514 6868 20402
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6000 19440 6052 19446
rect 6000 19382 6052 19388
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4712 18284 4764 18290
rect 4712 18226 4764 18232
rect 4724 17542 4752 18226
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 3595 16892 3903 16901
rect 3595 16890 3601 16892
rect 3657 16890 3681 16892
rect 3737 16890 3761 16892
rect 3817 16890 3841 16892
rect 3897 16890 3903 16892
rect 3657 16838 3659 16890
rect 3839 16838 3841 16890
rect 3595 16836 3601 16838
rect 3657 16836 3681 16838
rect 3737 16836 3761 16838
rect 3817 16836 3841 16838
rect 3897 16836 3903 16838
rect 3595 16827 3903 16836
rect 3516 16584 3568 16590
rect 3436 16544 3516 16572
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 3240 15700 3292 15706
rect 3160 15660 3240 15688
rect 2320 15642 2372 15648
rect 3240 15642 3292 15648
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2608 15094 2636 15302
rect 2596 15088 2648 15094
rect 2596 15030 2648 15036
rect 1492 15020 1544 15026
rect 1492 14962 1544 14968
rect 1504 14482 1532 14962
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 3068 13920 3096 15302
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 3160 14618 3188 14894
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3148 13932 3200 13938
rect 3068 13892 3148 13920
rect 3148 13874 3200 13880
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1596 11762 1624 12174
rect 2136 12164 2188 12170
rect 2136 12106 2188 12112
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1596 10130 1624 11698
rect 1780 11354 1808 11698
rect 2148 11354 2176 12106
rect 2884 11354 2912 12650
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 3068 11354 3096 11494
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2424 10810 2452 11086
rect 2792 10810 2820 11086
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2976 10606 3004 10950
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1596 9586 1624 10066
rect 1964 10062 1992 10406
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 2976 9722 3004 10542
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 3160 9654 3188 13874
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 992 8936 994 8945
rect 938 8871 994 8880
rect 1596 8498 1624 9522
rect 2240 9178 2268 9522
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1872 5030 1900 8910
rect 3252 6254 3280 15642
rect 3436 15434 3464 16544
rect 3516 16526 3568 16532
rect 4080 16522 4108 17002
rect 4448 16590 4476 17138
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3528 15706 3556 16390
rect 4255 16348 4563 16357
rect 4255 16346 4261 16348
rect 4317 16346 4341 16348
rect 4397 16346 4421 16348
rect 4477 16346 4501 16348
rect 4557 16346 4563 16348
rect 4317 16294 4319 16346
rect 4499 16294 4501 16346
rect 4255 16292 4261 16294
rect 4317 16292 4341 16294
rect 4397 16292 4421 16294
rect 4477 16292 4501 16294
rect 4557 16292 4563 16294
rect 4255 16283 4563 16292
rect 4632 16250 4660 16594
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 3595 15804 3903 15813
rect 3595 15802 3601 15804
rect 3657 15802 3681 15804
rect 3737 15802 3761 15804
rect 3817 15802 3841 15804
rect 3897 15802 3903 15804
rect 3657 15750 3659 15802
rect 3839 15750 3841 15802
rect 3595 15748 3601 15750
rect 3657 15748 3681 15750
rect 3737 15748 3761 15750
rect 3817 15748 3841 15750
rect 3897 15748 3903 15750
rect 3595 15739 3903 15748
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 4540 15570 4568 16050
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4632 15586 4660 15846
rect 4724 15706 4752 17138
rect 4908 16794 4936 18770
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5078 18456 5134 18465
rect 5078 18391 5134 18400
rect 5092 18358 5120 18391
rect 5080 18352 5132 18358
rect 5080 18294 5132 18300
rect 5552 18290 5580 18566
rect 5920 18426 5948 19314
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5920 18290 5948 18362
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5552 17678 5580 18226
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4816 16114 4844 16390
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5000 15706 5028 15846
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4528 15564 4580 15570
rect 4632 15558 4752 15586
rect 4528 15506 4580 15512
rect 3424 15428 3476 15434
rect 3424 15370 3476 15376
rect 3436 14890 3464 15370
rect 4080 15094 4108 15506
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4172 15162 4200 15302
rect 4255 15260 4563 15269
rect 4255 15258 4261 15260
rect 4317 15258 4341 15260
rect 4397 15258 4421 15260
rect 4477 15258 4501 15260
rect 4557 15258 4563 15260
rect 4317 15206 4319 15258
rect 4499 15206 4501 15258
rect 4255 15204 4261 15206
rect 4317 15204 4341 15206
rect 4397 15204 4421 15206
rect 4477 15204 4501 15206
rect 4557 15204 4563 15206
rect 4255 15195 4563 15204
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 3516 15088 3568 15094
rect 3516 15030 3568 15036
rect 4068 15088 4120 15094
rect 4120 15036 4292 15042
rect 4068 15030 4292 15036
rect 3424 14884 3476 14890
rect 3424 14826 3476 14832
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3344 14618 3372 14758
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3528 14414 3556 15030
rect 4080 15014 4292 15030
rect 4264 14958 4292 15014
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3595 14716 3903 14725
rect 3595 14714 3601 14716
rect 3657 14714 3681 14716
rect 3737 14714 3761 14716
rect 3817 14714 3841 14716
rect 3897 14714 3903 14716
rect 3657 14662 3659 14714
rect 3839 14662 3841 14714
rect 3595 14660 3601 14662
rect 3657 14660 3681 14662
rect 3737 14660 3761 14662
rect 3817 14660 3841 14662
rect 3897 14660 3903 14662
rect 3595 14651 3903 14660
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3988 14346 4016 14758
rect 4080 14618 4108 14894
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 3988 14074 4016 14282
rect 4172 14074 4200 14758
rect 4448 14618 4476 14962
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4540 14482 4568 14962
rect 4632 14958 4660 15438
rect 4724 15366 4752 15558
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4724 14890 4752 15302
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 4908 14618 4936 15302
rect 5000 15162 5028 15438
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 5092 14414 5120 14758
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 4255 14172 4563 14181
rect 4255 14170 4261 14172
rect 4317 14170 4341 14172
rect 4397 14170 4421 14172
rect 4477 14170 4501 14172
rect 4557 14170 4563 14172
rect 4317 14118 4319 14170
rect 4499 14118 4501 14170
rect 4255 14116 4261 14118
rect 4317 14116 4341 14118
rect 4397 14116 4421 14118
rect 4477 14116 4501 14118
rect 4557 14116 4563 14118
rect 4255 14107 4563 14116
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 5092 14006 5120 14350
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 5080 14000 5132 14006
rect 5080 13942 5132 13948
rect 3595 13628 3903 13637
rect 3595 13626 3601 13628
rect 3657 13626 3681 13628
rect 3737 13626 3761 13628
rect 3817 13626 3841 13628
rect 3897 13626 3903 13628
rect 3657 13574 3659 13626
rect 3839 13574 3841 13626
rect 3595 13572 3601 13574
rect 3657 13572 3681 13574
rect 3737 13572 3761 13574
rect 3817 13572 3841 13574
rect 3897 13572 3903 13574
rect 3595 13563 3903 13572
rect 4356 13394 4384 13942
rect 5184 13938 5212 17478
rect 5644 17320 5672 18158
rect 6012 18154 6040 19382
rect 6840 19378 6868 19450
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6104 18290 6132 18770
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 5552 17292 5672 17320
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 16114 5304 16934
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4356 13274 4384 13330
rect 4172 13246 4384 13274
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3528 12442 3556 12718
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 3595 12540 3903 12549
rect 3595 12538 3601 12540
rect 3657 12538 3681 12540
rect 3737 12538 3761 12540
rect 3817 12538 3841 12540
rect 3897 12538 3903 12540
rect 3657 12486 3659 12538
rect 3839 12486 3841 12538
rect 3595 12484 3601 12486
rect 3657 12484 3681 12486
rect 3737 12484 3761 12486
rect 3817 12484 3841 12486
rect 3897 12484 3903 12486
rect 3595 12475 3903 12484
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 4080 12374 4108 12650
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 3332 11620 3384 11626
rect 3332 11562 3384 11568
rect 3344 11132 3372 11562
rect 3436 11354 3464 12310
rect 4172 12238 4200 13246
rect 4255 13084 4563 13093
rect 4255 13082 4261 13084
rect 4317 13082 4341 13084
rect 4397 13082 4421 13084
rect 4477 13082 4501 13084
rect 4557 13082 4563 13084
rect 4317 13030 4319 13082
rect 4499 13030 4501 13082
rect 4255 13028 4261 13030
rect 4317 13028 4341 13030
rect 4397 13028 4421 13030
rect 4477 13028 4501 13030
rect 4557 13028 4563 13030
rect 4255 13019 4563 13028
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4448 12238 4476 12582
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 4172 11762 4200 12174
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4255 11996 4563 12005
rect 4255 11994 4261 11996
rect 4317 11994 4341 11996
rect 4397 11994 4421 11996
rect 4477 11994 4501 11996
rect 4557 11994 4563 11996
rect 4317 11942 4319 11994
rect 4499 11942 4501 11994
rect 4255 11940 4261 11942
rect 4317 11940 4341 11942
rect 4397 11940 4421 11942
rect 4477 11940 4501 11942
rect 4557 11940 4563 11942
rect 4255 11931 4563 11940
rect 4632 11898 4660 12038
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 3595 11452 3903 11461
rect 3595 11450 3601 11452
rect 3657 11450 3681 11452
rect 3737 11450 3761 11452
rect 3817 11450 3841 11452
rect 3897 11450 3903 11452
rect 3657 11398 3659 11450
rect 3839 11398 3841 11450
rect 3595 11396 3601 11398
rect 3657 11396 3681 11398
rect 3737 11396 3761 11398
rect 3817 11396 3841 11398
rect 3897 11396 3903 11398
rect 3595 11387 3903 11396
rect 3424 11348 3476 11354
rect 3476 11308 3556 11336
rect 3424 11290 3476 11296
rect 3528 11150 3556 11308
rect 4172 11218 4200 11698
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4264 11354 4292 11494
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 3424 11144 3476 11150
rect 3344 11104 3424 11132
rect 3424 11086 3476 11092
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3344 10674 3372 10950
rect 3896 10674 3924 10950
rect 4255 10908 4563 10917
rect 4255 10906 4261 10908
rect 4317 10906 4341 10908
rect 4397 10906 4421 10908
rect 4477 10906 4501 10908
rect 4557 10906 4563 10908
rect 4317 10854 4319 10906
rect 4499 10854 4501 10906
rect 4255 10852 4261 10854
rect 4317 10852 4341 10854
rect 4397 10852 4421 10854
rect 4477 10852 4501 10854
rect 4557 10852 4563 10854
rect 4255 10843 4563 10852
rect 4632 10674 4660 11154
rect 4908 11150 4936 12038
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 3344 10266 3372 10610
rect 3595 10364 3903 10373
rect 3595 10362 3601 10364
rect 3657 10362 3681 10364
rect 3737 10362 3761 10364
rect 3817 10362 3841 10364
rect 3897 10362 3903 10364
rect 3657 10310 3659 10362
rect 3839 10310 3841 10362
rect 3595 10308 3601 10310
rect 3657 10308 3681 10310
rect 3737 10308 3761 10310
rect 3817 10308 3841 10310
rect 3897 10308 3903 10310
rect 3595 10299 3903 10308
rect 5276 10266 5304 12174
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 4255 9820 4563 9829
rect 4255 9818 4261 9820
rect 4317 9818 4341 9820
rect 4397 9818 4421 9820
rect 4477 9818 4501 9820
rect 4557 9818 4563 9820
rect 4317 9766 4319 9818
rect 4499 9766 4501 9818
rect 4255 9764 4261 9766
rect 4317 9764 4341 9766
rect 4397 9764 4421 9766
rect 4477 9764 4501 9766
rect 4557 9764 4563 9766
rect 4255 9755 4563 9764
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3595 9276 3903 9285
rect 3595 9274 3601 9276
rect 3657 9274 3681 9276
rect 3737 9274 3761 9276
rect 3817 9274 3841 9276
rect 3897 9274 3903 9276
rect 3657 9222 3659 9274
rect 3839 9222 3841 9274
rect 3595 9220 3601 9222
rect 3657 9220 3681 9222
rect 3737 9220 3761 9222
rect 3817 9220 3841 9222
rect 3897 9220 3903 9222
rect 3595 9211 3903 9220
rect 3988 8634 4016 9318
rect 4080 9178 4108 9590
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4356 9178 4384 9454
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 5092 8974 5120 9318
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3528 7886 3556 8230
rect 3595 8188 3903 8197
rect 3595 8186 3601 8188
rect 3657 8186 3681 8188
rect 3737 8186 3761 8188
rect 3817 8186 3841 8188
rect 3897 8186 3903 8188
rect 3657 8134 3659 8186
rect 3839 8134 3841 8186
rect 3595 8132 3601 8134
rect 3657 8132 3681 8134
rect 3737 8132 3761 8134
rect 3817 8132 3841 8134
rect 3897 8132 3903 8134
rect 3595 8123 3903 8132
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3884 7880 3936 7886
rect 3936 7840 4016 7868
rect 3884 7822 3936 7828
rect 3988 7206 4016 7840
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3595 7100 3903 7109
rect 3595 7098 3601 7100
rect 3657 7098 3681 7100
rect 3737 7098 3761 7100
rect 3817 7098 3841 7100
rect 3897 7098 3903 7100
rect 3657 7046 3659 7098
rect 3839 7046 3841 7098
rect 3595 7044 3601 7046
rect 3657 7044 3681 7046
rect 3737 7044 3761 7046
rect 3817 7044 3841 7046
rect 3897 7044 3903 7046
rect 3595 7035 3903 7044
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3252 5914 3280 6190
rect 3595 6012 3903 6021
rect 3595 6010 3601 6012
rect 3657 6010 3681 6012
rect 3737 6010 3761 6012
rect 3817 6010 3841 6012
rect 3897 6010 3903 6012
rect 3657 5958 3659 6010
rect 3839 5958 3841 6010
rect 3595 5956 3601 5958
rect 3657 5956 3681 5958
rect 3737 5956 3761 5958
rect 3817 5956 3841 5958
rect 3897 5956 3903 5958
rect 3595 5947 3903 5956
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3988 5710 4016 7142
rect 4080 6798 4108 8910
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 7818 4200 8774
rect 4255 8732 4563 8741
rect 4255 8730 4261 8732
rect 4317 8730 4341 8732
rect 4397 8730 4421 8732
rect 4477 8730 4501 8732
rect 4557 8730 4563 8732
rect 4317 8678 4319 8730
rect 4499 8678 4501 8730
rect 4255 8676 4261 8678
rect 4317 8676 4341 8678
rect 4397 8676 4421 8678
rect 4477 8676 4501 8678
rect 4557 8676 4563 8678
rect 4255 8667 4563 8676
rect 5092 8294 5120 8910
rect 5276 8634 5304 9318
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 4255 7644 4563 7653
rect 4255 7642 4261 7644
rect 4317 7642 4341 7644
rect 4397 7642 4421 7644
rect 4477 7642 4501 7644
rect 4557 7642 4563 7644
rect 4317 7590 4319 7642
rect 4499 7590 4501 7642
rect 4255 7588 4261 7590
rect 4317 7588 4341 7590
rect 4397 7588 4421 7590
rect 4477 7588 4501 7590
rect 4557 7588 4563 7590
rect 4255 7579 4563 7588
rect 5092 7546 5120 8230
rect 5368 7886 5396 16050
rect 5552 16046 5580 17292
rect 6196 17270 6224 19314
rect 6276 19304 6328 19310
rect 6276 19246 6328 19252
rect 6288 18630 6316 19246
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6368 18692 6420 18698
rect 6368 18634 6420 18640
rect 6276 18624 6328 18630
rect 6276 18566 6328 18572
rect 6380 18426 6408 18634
rect 6368 18420 6420 18426
rect 6368 18362 6420 18368
rect 6564 18290 6592 19110
rect 6656 18698 6684 19110
rect 6736 18760 6788 18766
rect 6736 18702 6788 18708
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6656 18290 6684 18634
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6472 18170 6500 18226
rect 6748 18170 6776 18702
rect 6472 18142 6776 18170
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5644 16794 5672 17138
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5736 16250 5764 16458
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 6104 16114 6132 16934
rect 6472 16794 6500 18142
rect 6748 18086 6776 18142
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6368 16788 6420 16794
rect 6368 16730 6420 16736
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 6380 16114 6408 16730
rect 6564 16658 6592 17138
rect 6552 16652 6604 16658
rect 6472 16612 6552 16640
rect 6472 16114 6500 16612
rect 6552 16594 6604 16600
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 6564 15910 6592 16050
rect 6656 15978 6684 17138
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6564 15094 6592 15846
rect 6552 15088 6604 15094
rect 6552 15030 6604 15036
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5460 14074 5488 14418
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5644 14074 5672 14350
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5552 12442 5580 13874
rect 5828 13870 5856 14758
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 6012 13326 6040 14486
rect 6748 14414 6776 14962
rect 6840 14822 6868 19314
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7208 18834 7236 19110
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7300 18426 7328 20538
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 7668 19122 7696 20878
rect 7748 20868 7800 20874
rect 7748 20810 7800 20816
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 7760 20602 7788 20810
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 8680 20534 8708 20810
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 8668 20528 8720 20534
rect 8668 20470 8720 20476
rect 8885 20156 9193 20165
rect 8885 20154 8891 20156
rect 8947 20154 8971 20156
rect 9027 20154 9051 20156
rect 9107 20154 9131 20156
rect 9187 20154 9193 20156
rect 8947 20102 8949 20154
rect 9129 20102 9131 20154
rect 8885 20100 8891 20102
rect 8947 20100 8971 20102
rect 9027 20100 9051 20102
rect 9107 20100 9131 20102
rect 9187 20100 9193 20102
rect 8885 20091 9193 20100
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 7932 19168 7984 19174
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7116 16726 7144 17070
rect 7104 16720 7156 16726
rect 7104 16662 7156 16668
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6932 16250 6960 16526
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7116 16114 7144 16662
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7300 15706 7328 17138
rect 7392 16794 7420 18702
rect 7484 18290 7512 19110
rect 7668 19094 7788 19122
rect 7932 19110 7984 19116
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7484 16590 7512 16934
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7484 16114 7512 16390
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7484 15366 7512 16050
rect 7576 15502 7604 16934
rect 7668 16114 7696 18906
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7668 15502 7696 16050
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7668 15366 7696 15438
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 7024 14414 7052 14826
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7392 14498 7420 14758
rect 7484 14618 7512 15302
rect 7668 14890 7696 15302
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7392 14470 7512 14498
rect 7484 14414 7512 14470
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 6748 14074 6776 14350
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6932 13954 6960 14282
rect 6656 13938 6960 13954
rect 7024 13938 7052 14350
rect 6644 13932 6960 13938
rect 6696 13926 6960 13932
rect 6644 13874 6696 13880
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 6840 12918 6868 13806
rect 6932 13190 6960 13926
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7024 13818 7052 13874
rect 7024 13790 7144 13818
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6932 12850 6960 13126
rect 7024 12986 7052 13670
rect 7116 13530 7144 13790
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7116 12850 7144 13466
rect 7392 12986 7420 13874
rect 7484 13258 7512 14350
rect 7760 14278 7788 19094
rect 7944 18766 7972 19110
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 8312 18698 8340 19110
rect 8404 18834 8432 19246
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8220 18290 8248 18566
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7852 15706 7880 17138
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8220 16726 8248 17002
rect 8496 16998 8524 18158
rect 8588 18154 8616 19450
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 8668 19236 8720 19242
rect 8668 19178 8720 19184
rect 8680 18698 8708 19178
rect 8885 19068 9193 19077
rect 8885 19066 8891 19068
rect 8947 19066 8971 19068
rect 9027 19066 9051 19068
rect 9107 19066 9131 19068
rect 9187 19066 9193 19068
rect 8947 19014 8949 19066
rect 9129 19014 9131 19066
rect 8885 19012 8891 19014
rect 8947 19012 8971 19014
rect 9027 19012 9051 19014
rect 9107 19012 9131 19014
rect 9187 19012 9193 19014
rect 8885 19003 9193 19012
rect 9232 18970 9260 19314
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8864 18426 8892 18770
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 9232 18154 9260 18634
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 8220 16114 8248 16662
rect 8496 16522 8524 16934
rect 8484 16516 8536 16522
rect 8484 16458 8536 16464
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7852 13326 7880 14418
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8036 14074 8064 14350
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8312 13938 8340 16186
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8404 15026 8432 15506
rect 8496 15094 8524 16458
rect 8588 16454 8616 17070
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 8588 15638 8616 16390
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 8484 15088 8536 15094
rect 8484 15030 8536 15036
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8496 14618 8524 15030
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8496 14498 8524 14554
rect 8772 14550 8800 18022
rect 8885 17980 9193 17989
rect 8885 17978 8891 17980
rect 8947 17978 8971 17980
rect 9027 17978 9051 17980
rect 9107 17978 9131 17980
rect 9187 17978 9193 17980
rect 8947 17926 8949 17978
rect 9129 17926 9131 17978
rect 8885 17924 8891 17926
rect 8947 17924 8971 17926
rect 9027 17924 9051 17926
rect 9107 17924 9131 17926
rect 9187 17924 9193 17926
rect 8885 17915 9193 17924
rect 9324 17678 9352 20742
rect 9545 20700 9853 20709
rect 9545 20698 9551 20700
rect 9607 20698 9631 20700
rect 9687 20698 9711 20700
rect 9767 20698 9791 20700
rect 9847 20698 9853 20700
rect 9607 20646 9609 20698
rect 9789 20646 9791 20698
rect 9545 20644 9551 20646
rect 9607 20644 9631 20646
rect 9687 20644 9711 20646
rect 9767 20644 9791 20646
rect 9847 20644 9853 20646
rect 9545 20635 9853 20644
rect 9545 19612 9853 19621
rect 9545 19610 9551 19612
rect 9607 19610 9631 19612
rect 9687 19610 9711 19612
rect 9767 19610 9791 19612
rect 9847 19610 9853 19612
rect 9607 19558 9609 19610
rect 9789 19558 9791 19610
rect 9545 19556 9551 19558
rect 9607 19556 9631 19558
rect 9687 19556 9711 19558
rect 9767 19556 9791 19558
rect 9847 19556 9853 19558
rect 9545 19547 9853 19556
rect 9968 18766 9996 20896
rect 10232 20868 10284 20874
rect 10232 20810 10284 20816
rect 10244 20602 10272 20810
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10336 19360 10364 20742
rect 10428 20466 10456 21082
rect 10796 20942 10824 21286
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10796 20602 10824 20878
rect 10980 20806 11008 21490
rect 11992 21146 12020 21678
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 11980 21140 12032 21146
rect 12032 21100 12112 21128
rect 11980 21082 12032 21088
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 11164 20482 11192 20742
rect 10980 20466 11192 20482
rect 11256 20466 11284 20742
rect 11336 20528 11388 20534
rect 11336 20470 11388 20476
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10968 20460 11192 20466
rect 11020 20454 11192 20460
rect 10968 20402 11020 20408
rect 11164 20262 11192 20454
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11164 19378 11192 20198
rect 11348 19417 11376 20470
rect 12084 20466 12112 21100
rect 12176 20602 12204 21898
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12268 20602 12296 21082
rect 12164 20596 12216 20602
rect 12164 20538 12216 20544
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 12360 20466 12388 21898
rect 12728 21146 12756 22034
rect 13004 21146 13032 22102
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 13096 21690 13124 21966
rect 13464 21690 13492 22578
rect 13544 22568 13596 22574
rect 13544 22510 13596 22516
rect 13084 21684 13136 21690
rect 13084 21626 13136 21632
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13096 21146 13124 21626
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 12256 20324 12308 20330
rect 12256 20266 12308 20272
rect 11334 19408 11390 19417
rect 10416 19372 10468 19378
rect 10336 19332 10416 19360
rect 10416 19314 10468 19320
rect 11152 19372 11204 19378
rect 12162 19408 12218 19417
rect 11334 19343 11390 19352
rect 11888 19372 11940 19378
rect 11152 19314 11204 19320
rect 12162 19343 12218 19352
rect 11888 19314 11940 19320
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10244 18766 10272 19110
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 9545 18524 9853 18533
rect 9545 18522 9551 18524
rect 9607 18522 9631 18524
rect 9687 18522 9711 18524
rect 9767 18522 9791 18524
rect 9847 18522 9853 18524
rect 9607 18470 9609 18522
rect 9789 18470 9791 18522
rect 9545 18468 9551 18470
rect 9607 18468 9631 18470
rect 9687 18468 9711 18470
rect 9767 18468 9791 18470
rect 9847 18468 9853 18470
rect 9545 18459 9853 18468
rect 9680 18216 9732 18222
rect 9968 18204 9996 18702
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 10244 18290 10272 18566
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 9732 18176 9996 18204
rect 9680 18158 9732 18164
rect 9312 17672 9364 17678
rect 9232 17632 9312 17660
rect 9232 17241 9260 17632
rect 9312 17614 9364 17620
rect 9312 17536 9364 17542
rect 9692 17524 9720 18158
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 9312 17478 9364 17484
rect 9416 17496 9720 17524
rect 9218 17232 9274 17241
rect 9324 17202 9352 17478
rect 9218 17167 9274 17176
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9416 16998 9444 17496
rect 9545 17436 9853 17445
rect 9545 17434 9551 17436
rect 9607 17434 9631 17436
rect 9687 17434 9711 17436
rect 9767 17434 9791 17436
rect 9847 17434 9853 17436
rect 9607 17382 9609 17434
rect 9789 17382 9791 17434
rect 9545 17380 9551 17382
rect 9607 17380 9631 17382
rect 9687 17380 9711 17382
rect 9767 17380 9791 17382
rect 9847 17380 9853 17382
rect 9545 17371 9853 17380
rect 9496 17264 9548 17270
rect 9494 17232 9496 17241
rect 9548 17232 9550 17241
rect 9494 17167 9550 17176
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 8885 16892 9193 16901
rect 8885 16890 8891 16892
rect 8947 16890 8971 16892
rect 9027 16890 9051 16892
rect 9107 16890 9131 16892
rect 9187 16890 9193 16892
rect 8947 16838 8949 16890
rect 9129 16838 9131 16890
rect 8885 16836 8891 16838
rect 8947 16836 8971 16838
rect 9027 16836 9051 16838
rect 9107 16836 9131 16838
rect 9187 16836 9193 16838
rect 8885 16827 9193 16836
rect 9416 16658 9444 16934
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9416 16250 9444 16594
rect 9508 16590 9536 17167
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9772 16584 9824 16590
rect 9968 16572 9996 17818
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 10060 16998 10088 17614
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 9824 16544 9996 16572
rect 9772 16526 9824 16532
rect 9545 16348 9853 16357
rect 9545 16346 9551 16348
rect 9607 16346 9631 16348
rect 9687 16346 9711 16348
rect 9767 16346 9791 16348
rect 9847 16346 9853 16348
rect 9607 16294 9609 16346
rect 9789 16294 9791 16346
rect 9545 16292 9551 16294
rect 9607 16292 9631 16294
rect 9687 16292 9711 16294
rect 9767 16292 9791 16294
rect 9847 16292 9853 16294
rect 9545 16283 9853 16292
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 8885 15804 9193 15813
rect 8885 15802 8891 15804
rect 8947 15802 8971 15804
rect 9027 15802 9051 15804
rect 9107 15802 9131 15804
rect 9187 15802 9193 15804
rect 8947 15750 8949 15802
rect 9129 15750 9131 15802
rect 8885 15748 8891 15750
rect 8947 15748 8971 15750
rect 9027 15748 9051 15750
rect 9107 15748 9131 15750
rect 9187 15748 9193 15750
rect 8885 15739 9193 15748
rect 9232 15570 9260 16050
rect 10152 15910 10180 17478
rect 10336 17338 10364 17546
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9545 15260 9853 15269
rect 9545 15258 9551 15260
rect 9607 15258 9631 15260
rect 9687 15258 9711 15260
rect 9767 15258 9791 15260
rect 9847 15258 9853 15260
rect 9607 15206 9609 15258
rect 9789 15206 9791 15258
rect 9545 15204 9551 15206
rect 9607 15204 9631 15206
rect 9687 15204 9711 15206
rect 9767 15204 9791 15206
rect 9847 15204 9853 15206
rect 9545 15195 9853 15204
rect 8885 14716 9193 14725
rect 8885 14714 8891 14716
rect 8947 14714 8971 14716
rect 9027 14714 9051 14716
rect 9107 14714 9131 14716
rect 9187 14714 9193 14716
rect 8947 14662 8949 14714
rect 9129 14662 9131 14714
rect 8885 14660 8891 14662
rect 8947 14660 8971 14662
rect 9027 14660 9051 14662
rect 9107 14660 9131 14662
rect 9187 14660 9193 14662
rect 8885 14651 9193 14660
rect 8404 14470 8524 14498
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 8404 14414 8432 14470
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8404 13938 8432 14214
rect 8496 14074 8524 14214
rect 8680 14074 8708 14486
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5552 11898 5580 12174
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5736 10470 5764 12174
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10062 5764 10406
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5552 9042 5580 9522
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5644 9178 5672 9318
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5356 7880 5408 7886
rect 5276 7840 5356 7868
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5184 7410 5212 7686
rect 5276 7478 5304 7840
rect 5356 7822 5408 7828
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4080 6458 4108 6734
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4172 6458 4200 6598
rect 4255 6556 4563 6565
rect 4255 6554 4261 6556
rect 4317 6554 4341 6556
rect 4397 6554 4421 6556
rect 4477 6554 4501 6556
rect 4557 6554 4563 6556
rect 4317 6502 4319 6554
rect 4499 6502 4501 6554
rect 4255 6500 4261 6502
rect 4317 6500 4341 6502
rect 4397 6500 4421 6502
rect 4477 6500 4501 6502
rect 4557 6500 4563 6502
rect 4255 6491 4563 6500
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4908 6390 4936 6598
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 3595 4924 3903 4933
rect 3595 4922 3601 4924
rect 3657 4922 3681 4924
rect 3737 4922 3761 4924
rect 3817 4922 3841 4924
rect 3897 4922 3903 4924
rect 3657 4870 3659 4922
rect 3839 4870 3841 4922
rect 3595 4868 3601 4870
rect 3657 4868 3681 4870
rect 3737 4868 3761 4870
rect 3817 4868 3841 4870
rect 3897 4868 3903 4870
rect 3595 4859 3903 4868
rect 3595 3836 3903 3845
rect 3595 3834 3601 3836
rect 3657 3834 3681 3836
rect 3737 3834 3761 3836
rect 3817 3834 3841 3836
rect 3897 3834 3903 3836
rect 3657 3782 3659 3834
rect 3839 3782 3841 3834
rect 3595 3780 3601 3782
rect 3657 3780 3681 3782
rect 3737 3780 3761 3782
rect 3817 3780 3841 3782
rect 3897 3780 3903 3782
rect 3595 3771 3903 3780
rect 4172 3058 4200 5646
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4255 5468 4563 5477
rect 4255 5466 4261 5468
rect 4317 5466 4341 5468
rect 4397 5466 4421 5468
rect 4477 5466 4501 5468
rect 4557 5466 4563 5468
rect 4317 5414 4319 5466
rect 4499 5414 4501 5466
rect 4255 5412 4261 5414
rect 4317 5412 4341 5414
rect 4397 5412 4421 5414
rect 4477 5412 4501 5414
rect 4557 5412 4563 5414
rect 4255 5403 4563 5412
rect 4632 5370 4660 5578
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4908 5234 4936 6326
rect 5552 6254 5580 7686
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5736 6730 5764 7142
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5552 5778 5580 6190
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 5092 4622 5120 5170
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4255 4380 4563 4389
rect 4255 4378 4261 4380
rect 4317 4378 4341 4380
rect 4397 4378 4421 4380
rect 4477 4378 4501 4380
rect 4557 4378 4563 4380
rect 4317 4326 4319 4378
rect 4499 4326 4501 4378
rect 4255 4324 4261 4326
rect 4317 4324 4341 4326
rect 4397 4324 4421 4326
rect 4477 4324 4501 4326
rect 4557 4324 4563 4326
rect 4255 4315 4563 4324
rect 4816 4078 4844 4558
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 4146 5396 4490
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4255 3292 4563 3301
rect 4255 3290 4261 3292
rect 4317 3290 4341 3292
rect 4397 3290 4421 3292
rect 4477 3290 4501 3292
rect 4557 3290 4563 3292
rect 4317 3238 4319 3290
rect 4499 3238 4501 3290
rect 4255 3236 4261 3238
rect 4317 3236 4341 3238
rect 4397 3236 4421 3238
rect 4477 3236 4501 3238
rect 4557 3236 4563 3238
rect 4255 3227 4563 3236
rect 4632 3194 4660 3878
rect 5092 3466 5120 3878
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 5184 3194 5212 4082
rect 5552 3534 5580 5714
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5644 5234 5672 5510
rect 5828 5234 5856 12378
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 10606 5948 11494
rect 6012 10742 6040 12038
rect 8680 11898 8708 12038
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6196 11014 6224 11630
rect 6380 11286 6408 11766
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6564 11354 6592 11494
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6380 10810 6408 11086
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5920 10130 5948 10542
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 6380 9994 6408 10746
rect 6564 10674 6592 10950
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6564 9994 6592 10610
rect 6656 10470 6684 11222
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6748 10266 6776 11766
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6840 10538 6868 11154
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7024 10674 7052 10950
rect 7116 10810 7144 11698
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7300 10810 7328 11494
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7760 10810 7788 11018
rect 8036 10810 8064 11698
rect 8772 11286 8800 14486
rect 9232 13734 9260 14486
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 8885 13628 9193 13637
rect 8885 13626 8891 13628
rect 8947 13626 8971 13628
rect 9027 13626 9051 13628
rect 9107 13626 9131 13628
rect 9187 13626 9193 13628
rect 8947 13574 8949 13626
rect 9129 13574 9131 13626
rect 8885 13572 8891 13574
rect 8947 13572 8971 13574
rect 9027 13572 9051 13574
rect 9107 13572 9131 13574
rect 9187 13572 9193 13574
rect 8885 13563 9193 13572
rect 9232 13394 9260 13670
rect 9324 13462 9352 14282
rect 9508 14260 9536 14350
rect 9416 14232 9536 14260
rect 10048 14272 10100 14278
rect 9416 13530 9444 14232
rect 10048 14214 10100 14220
rect 9545 14172 9853 14181
rect 9545 14170 9551 14172
rect 9607 14170 9631 14172
rect 9687 14170 9711 14172
rect 9767 14170 9791 14172
rect 9847 14170 9853 14172
rect 9607 14118 9609 14170
rect 9789 14118 9791 14170
rect 9545 14116 9551 14118
rect 9607 14116 9631 14118
rect 9687 14116 9711 14118
rect 9767 14116 9791 14118
rect 9847 14116 9853 14118
rect 9545 14107 9853 14116
rect 10060 13938 10088 14214
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 10152 13326 10180 14350
rect 10244 14074 10272 14350
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10244 13802 10272 14010
rect 10232 13796 10284 13802
rect 10232 13738 10284 13744
rect 10244 13394 10272 13738
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 9545 13084 9853 13093
rect 9545 13082 9551 13084
rect 9607 13082 9631 13084
rect 9687 13082 9711 13084
rect 9767 13082 9791 13084
rect 9847 13082 9853 13084
rect 9607 13030 9609 13082
rect 9789 13030 9791 13082
rect 9545 13028 9551 13030
rect 9607 13028 9631 13030
rect 9687 13028 9711 13030
rect 9767 13028 9791 13030
rect 9847 13028 9853 13030
rect 9545 13019 9853 13028
rect 8885 12540 9193 12549
rect 8885 12538 8891 12540
rect 8947 12538 8971 12540
rect 9027 12538 9051 12540
rect 9107 12538 9131 12540
rect 9187 12538 9193 12540
rect 8947 12486 8949 12538
rect 9129 12486 9131 12538
rect 8885 12484 8891 12486
rect 8947 12484 8971 12486
rect 9027 12484 9051 12486
rect 9107 12484 9131 12486
rect 9187 12484 9193 12486
rect 8885 12475 9193 12484
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9545 11996 9853 12005
rect 9545 11994 9551 11996
rect 9607 11994 9631 11996
rect 9687 11994 9711 11996
rect 9767 11994 9791 11996
rect 9847 11994 9853 11996
rect 9607 11942 9609 11994
rect 9789 11942 9791 11994
rect 9545 11940 9551 11942
rect 9607 11940 9631 11942
rect 9687 11940 9711 11942
rect 9767 11940 9791 11942
rect 9847 11940 9853 11942
rect 9545 11931 9853 11940
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 8885 11452 9193 11461
rect 8885 11450 8891 11452
rect 8947 11450 8971 11452
rect 9027 11450 9051 11452
rect 9107 11450 9131 11452
rect 9187 11450 9193 11452
rect 8947 11398 8949 11450
rect 9129 11398 9131 11450
rect 8885 11396 8891 11398
rect 8947 11396 8971 11398
rect 9027 11396 9051 11398
rect 9107 11396 9131 11398
rect 9187 11396 9193 11398
rect 8885 11387 9193 11396
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6828 10532 6880 10538
rect 6828 10474 6880 10480
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6104 9178 6132 9318
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6104 8634 6132 8910
rect 6380 8634 6408 9522
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7300 8838 7328 9386
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6104 8022 6132 8570
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6104 7546 6132 7958
rect 6932 7954 6960 8366
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6840 7478 6868 7754
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6932 7410 6960 7686
rect 7024 7546 7052 8502
rect 7392 8498 7420 9318
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7116 7546 7144 7822
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7392 7410 7420 8434
rect 7668 8090 7696 8434
rect 7760 8090 7788 9522
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8128 9178 8156 9318
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8220 8974 8248 9318
rect 8312 9178 8340 9522
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7484 7410 7512 7958
rect 7852 7954 7880 8366
rect 8036 7954 8064 8774
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5644 4078 5672 4422
rect 5920 4078 5948 4626
rect 6104 4622 6132 5170
rect 6288 4826 6316 5782
rect 6472 5642 6500 6666
rect 7208 6458 7236 6802
rect 7300 6798 7328 7346
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7300 6458 7328 6734
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5710 6960 6190
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6932 5302 6960 5646
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 7116 5234 7144 6258
rect 7300 5846 7328 6394
rect 7392 6254 7420 7346
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 5920 2922 5948 4014
rect 6104 3194 6132 4558
rect 6288 3194 6316 4762
rect 7392 4622 7420 6054
rect 7576 5914 7604 6258
rect 7852 6254 7880 7890
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 8036 7002 8064 7754
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 8036 6798 8064 6938
rect 8220 6882 8248 8910
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8312 7342 8340 8434
rect 8404 8362 8432 9318
rect 8680 8838 8708 9454
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8430 8708 8774
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8404 7410 8432 8298
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8220 6854 8340 6882
rect 8496 6866 8524 8298
rect 8772 7750 8800 11222
rect 9692 11098 9720 11834
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9784 11354 9812 11630
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9968 11150 9996 12174
rect 10152 11830 10180 13262
rect 10336 12288 10364 16050
rect 10428 12442 10456 19314
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10888 18970 10916 19110
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10888 18290 10916 18906
rect 11164 18630 11192 19314
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11256 18426 11284 18634
rect 11532 18426 11560 18702
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11348 17882 11376 18226
rect 11336 17876 11388 17882
rect 11336 17818 11388 17824
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11256 16726 11284 17070
rect 11348 16998 11376 17614
rect 11336 16992 11388 16998
rect 11612 16992 11664 16998
rect 11388 16952 11560 16980
rect 11336 16934 11388 16940
rect 11244 16720 11296 16726
rect 11244 16662 11296 16668
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 11348 16046 11376 16526
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11440 16182 11468 16390
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 11532 16114 11560 16952
rect 11612 16934 11664 16940
rect 11624 16182 11652 16934
rect 11612 16176 11664 16182
rect 11612 16118 11664 16124
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10888 14074 10916 14214
rect 10980 14074 11008 14350
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10520 12442 10548 13330
rect 10796 13258 10824 13874
rect 11348 13870 11376 15982
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11624 13870 11652 14214
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10244 12260 10364 12288
rect 10244 11898 10272 12260
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10336 11898 10364 12106
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 10244 11370 10272 11834
rect 10428 11626 10456 12378
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 10796 11762 10824 12038
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10244 11342 10456 11370
rect 10612 11354 10640 11494
rect 9600 11082 9720 11098
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9588 11076 9720 11082
rect 9640 11070 9720 11076
rect 9588 11018 9640 11024
rect 9545 10908 9853 10917
rect 9545 10906 9551 10908
rect 9607 10906 9631 10908
rect 9687 10906 9711 10908
rect 9767 10906 9791 10908
rect 9847 10906 9853 10908
rect 9607 10854 9609 10906
rect 9789 10854 9791 10906
rect 9545 10852 9551 10854
rect 9607 10852 9631 10854
rect 9687 10852 9711 10854
rect 9767 10852 9791 10854
rect 9847 10852 9853 10854
rect 9545 10843 9853 10852
rect 9968 10606 9996 11086
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10152 10810 10180 10950
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 8885 10364 9193 10373
rect 8885 10362 8891 10364
rect 8947 10362 8971 10364
rect 9027 10362 9051 10364
rect 9107 10362 9131 10364
rect 9187 10362 9193 10364
rect 8947 10310 8949 10362
rect 9129 10310 9131 10362
rect 8885 10308 8891 10310
rect 8947 10308 8971 10310
rect 9027 10308 9051 10310
rect 9107 10308 9131 10310
rect 9187 10308 9193 10310
rect 8885 10299 9193 10308
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9324 9654 9352 9862
rect 9545 9820 9853 9829
rect 9545 9818 9551 9820
rect 9607 9818 9631 9820
rect 9687 9818 9711 9820
rect 9767 9818 9791 9820
rect 9847 9818 9853 9820
rect 9607 9766 9609 9818
rect 9789 9766 9791 9818
rect 9545 9764 9551 9766
rect 9607 9764 9631 9766
rect 9687 9764 9711 9766
rect 9767 9764 9791 9766
rect 9847 9764 9853 9766
rect 9545 9755 9853 9764
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9968 9518 9996 10542
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10060 9722 10088 9998
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 8885 9276 9193 9285
rect 8885 9274 8891 9276
rect 8947 9274 8971 9276
rect 9027 9274 9051 9276
rect 9107 9274 9131 9276
rect 9187 9274 9193 9276
rect 8947 9222 8949 9274
rect 9129 9222 9131 9274
rect 8885 9220 8891 9222
rect 8947 9220 8971 9222
rect 9027 9220 9051 9222
rect 9107 9220 9131 9222
rect 9187 9220 9193 9222
rect 8885 9211 9193 9220
rect 10060 9178 10088 9454
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9048 8634 9076 8978
rect 9220 8968 9272 8974
rect 9272 8928 9444 8956
rect 9220 8910 9272 8916
rect 9416 8922 9444 8928
rect 9416 8906 9536 8922
rect 9416 8900 9548 8906
rect 9416 8894 9496 8900
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9140 8566 9168 8774
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 8885 8188 9193 8197
rect 8885 8186 8891 8188
rect 8947 8186 8971 8188
rect 9027 8186 9051 8188
rect 9107 8186 9131 8188
rect 9187 8186 9193 8188
rect 8947 8134 8949 8186
rect 9129 8134 9131 8186
rect 8885 8132 8891 8134
rect 8947 8132 8971 8134
rect 9027 8132 9051 8134
rect 9107 8132 9131 8134
rect 9187 8132 9193 8134
rect 8885 8123 9193 8132
rect 9232 8090 9260 8434
rect 9324 8294 9352 8774
rect 9416 8634 9444 8894
rect 9496 8842 9548 8848
rect 9545 8732 9853 8741
rect 9545 8730 9551 8732
rect 9607 8730 9631 8732
rect 9687 8730 9711 8732
rect 9767 8730 9791 8732
rect 9847 8730 9853 8732
rect 9607 8678 9609 8730
rect 9789 8678 9791 8730
rect 9545 8676 9551 8678
rect 9607 8676 9631 8678
rect 9687 8676 9711 8678
rect 9767 8676 9791 8678
rect 9847 8676 9853 8678
rect 9545 8667 9853 8676
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9864 8560 9916 8566
rect 9862 8528 9864 8537
rect 9916 8528 9918 8537
rect 9588 8492 9640 8498
rect 9862 8463 9918 8472
rect 9588 8434 9640 8440
rect 9600 8362 9628 8434
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8885 7100 9193 7109
rect 8885 7098 8891 7100
rect 8947 7098 8971 7100
rect 9027 7098 9051 7100
rect 9107 7098 9131 7100
rect 9187 7098 9193 7100
rect 8947 7046 8949 7098
rect 9129 7046 9131 7098
rect 8885 7044 8891 7046
rect 8947 7044 8971 7046
rect 9027 7044 9051 7046
rect 9107 7044 9131 7046
rect 9187 7044 9193 7046
rect 8885 7035 9193 7044
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8024 6384 8076 6390
rect 8024 6326 8076 6332
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7576 5370 7604 5850
rect 8036 5642 8064 6326
rect 8220 6254 8248 6666
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8312 6186 8340 6854
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 9416 6798 9444 8298
rect 9600 8022 9628 8298
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9876 7750 9904 8463
rect 9968 7954 9996 8570
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 10060 7886 10088 9114
rect 10152 8838 10180 9522
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10244 8974 10272 9454
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10152 7886 10180 8774
rect 10244 8537 10272 8910
rect 10230 8528 10286 8537
rect 10230 8463 10286 8472
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10244 7886 10272 8230
rect 10336 8090 10364 9998
rect 10428 9586 10456 11342
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10784 9648 10836 9654
rect 10888 9602 10916 11834
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10836 9596 10916 9602
rect 10784 9590 10916 9596
rect 10416 9580 10468 9586
rect 10600 9580 10652 9586
rect 10468 9540 10548 9568
rect 10416 9522 10468 9528
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10428 9178 10456 9386
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10520 9110 10548 9540
rect 10600 9522 10652 9528
rect 10796 9574 10916 9590
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10428 8498 10456 8978
rect 10520 8974 10548 9046
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10612 8634 10640 9522
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8634 10732 8774
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10796 8514 10824 9574
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10520 8486 10824 8514
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 9864 7744 9916 7750
rect 9916 7692 9996 7698
rect 9864 7686 9996 7692
rect 9876 7670 9996 7686
rect 9545 7644 9853 7653
rect 9545 7642 9551 7644
rect 9607 7642 9631 7644
rect 9687 7642 9711 7644
rect 9767 7642 9791 7644
rect 9847 7642 9853 7644
rect 9607 7590 9609 7642
rect 9789 7590 9791 7642
rect 9545 7588 9551 7590
rect 9607 7588 9631 7590
rect 9687 7588 9711 7590
rect 9767 7588 9791 7590
rect 9847 7588 9853 7590
rect 9545 7579 9853 7588
rect 9864 6860 9916 6866
rect 9968 6848 9996 7670
rect 10336 7206 10364 7890
rect 10428 7886 10456 8230
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 9916 6820 9996 6848
rect 9864 6802 9916 6808
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 6458 8432 6598
rect 8588 6458 8616 6734
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8312 5710 8340 6122
rect 8588 5914 8616 6394
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8680 5710 8708 6598
rect 9232 6458 9260 6734
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 8772 5794 8800 6258
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 8885 6012 9193 6021
rect 8885 6010 8891 6012
rect 8947 6010 8971 6012
rect 9027 6010 9051 6012
rect 9107 6010 9131 6012
rect 9187 6010 9193 6012
rect 8947 5958 8949 6010
rect 9129 5958 9131 6010
rect 8885 5956 8891 5958
rect 8947 5956 8971 5958
rect 9027 5956 9051 5958
rect 9107 5956 9131 5958
rect 9187 5956 9193 5958
rect 8885 5947 9193 5956
rect 8772 5766 8892 5794
rect 9232 5778 9260 6190
rect 8864 5710 8892 5766
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 4758 7512 5170
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7576 4826 7604 4966
rect 7668 4826 7696 4966
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7760 4758 7788 5102
rect 7472 4752 7524 4758
rect 7748 4752 7800 4758
rect 7524 4700 7696 4706
rect 7472 4694 7696 4700
rect 7748 4694 7800 4700
rect 7484 4690 7696 4694
rect 7484 4684 7708 4690
rect 7484 4678 7656 4684
rect 7656 4626 7708 4632
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6840 3466 6868 3878
rect 6932 3670 6960 3878
rect 7300 3738 7328 4558
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6840 3194 6868 3402
rect 6932 3194 6960 3606
rect 7944 3534 7972 4150
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8036 3670 8064 4082
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6288 2922 6592 2938
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 6276 2916 6592 2922
rect 6328 2910 6592 2916
rect 6276 2858 6328 2864
rect 6564 2854 6592 2910
rect 8036 2854 8064 3606
rect 8128 3534 8156 4422
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8220 3194 8248 3878
rect 8312 3194 8340 5646
rect 9324 5642 9352 6258
rect 9416 5914 9444 6734
rect 9864 6724 9916 6730
rect 9916 6684 9996 6712
rect 9864 6666 9916 6672
rect 9545 6556 9853 6565
rect 9545 6554 9551 6556
rect 9607 6554 9631 6556
rect 9687 6554 9711 6556
rect 9767 6554 9791 6556
rect 9847 6554 9853 6556
rect 9607 6502 9609 6554
rect 9789 6502 9791 6554
rect 9545 6500 9551 6502
rect 9607 6500 9631 6502
rect 9687 6500 9711 6502
rect 9767 6500 9791 6502
rect 9847 6500 9853 6502
rect 9545 6491 9853 6500
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9600 6118 9628 6190
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 4146 8708 5510
rect 8885 4924 9193 4933
rect 8885 4922 8891 4924
rect 8947 4922 8971 4924
rect 9027 4922 9051 4924
rect 9107 4922 9131 4924
rect 9187 4922 9193 4924
rect 8947 4870 8949 4922
rect 9129 4870 9131 4922
rect 8885 4868 8891 4870
rect 8947 4868 8971 4870
rect 9027 4868 9051 4870
rect 9107 4868 9131 4870
rect 9187 4868 9193 4870
rect 8885 4859 9193 4868
rect 9232 4146 9260 5578
rect 9324 5234 9352 5578
rect 9416 5574 9444 5850
rect 9784 5692 9812 5850
rect 9876 5794 9904 6190
rect 9968 5914 9996 6684
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10060 6458 10088 6598
rect 10428 6458 10456 6734
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9876 5766 9996 5794
rect 9864 5704 9916 5710
rect 9678 5672 9734 5681
rect 9784 5664 9864 5692
rect 9864 5646 9916 5652
rect 9678 5607 9680 5616
rect 9732 5607 9734 5616
rect 9680 5578 9732 5584
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9545 5468 9853 5477
rect 9545 5466 9551 5468
rect 9607 5466 9631 5468
rect 9687 5466 9711 5468
rect 9767 5466 9791 5468
rect 9847 5466 9853 5468
rect 9607 5414 9609 5466
rect 9789 5414 9791 5466
rect 9545 5412 9551 5414
rect 9607 5412 9631 5414
rect 9687 5412 9711 5414
rect 9767 5412 9791 5414
rect 9847 5412 9853 5414
rect 9545 5403 9853 5412
rect 9968 5386 9996 5766
rect 9876 5358 9996 5386
rect 9876 5234 9904 5358
rect 10060 5234 10088 6394
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9545 4380 9853 4389
rect 9545 4378 9551 4380
rect 9607 4378 9631 4380
rect 9687 4378 9711 4380
rect 9767 4378 9791 4380
rect 9847 4378 9853 4380
rect 9607 4326 9609 4378
rect 9789 4326 9791 4378
rect 9545 4324 9551 4326
rect 9607 4324 9631 4326
rect 9687 4324 9711 4326
rect 9767 4324 9791 4326
rect 9847 4324 9853 4326
rect 9545 4315 9853 4324
rect 9772 4208 9824 4214
rect 9770 4176 9772 4185
rect 9824 4176 9826 4185
rect 9416 4146 9628 4162
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9416 4140 9640 4146
rect 9416 4134 9588 4140
rect 8404 3738 8432 4082
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8496 3534 8524 3878
rect 8680 3602 8708 4082
rect 8885 3836 9193 3845
rect 8885 3834 8891 3836
rect 8947 3834 8971 3836
rect 9027 3834 9051 3836
rect 9107 3834 9131 3836
rect 9187 3834 9193 3836
rect 8947 3782 8949 3834
rect 9129 3782 9131 3834
rect 8885 3780 8891 3782
rect 8947 3780 8971 3782
rect 9027 3780 9051 3782
rect 9107 3780 9131 3782
rect 9187 3780 9193 3782
rect 8885 3771 9193 3780
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 9232 3534 9260 4082
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8496 3058 8524 3334
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 9232 2854 9260 3470
rect 9416 3398 9444 4134
rect 9770 4111 9826 4120
rect 9588 4082 9640 4088
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9600 3670 9628 3946
rect 9784 3738 9812 4014
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9588 3664 9640 3670
rect 9588 3606 9640 3612
rect 10428 3398 10456 5646
rect 10520 3534 10548 8486
rect 10692 8424 10744 8430
rect 10744 8372 10916 8378
rect 10692 8366 10916 8372
rect 10704 8350 10916 8366
rect 10888 8106 10916 8350
rect 10980 8294 11008 11086
rect 11164 11082 11192 11494
rect 11256 11082 11284 12038
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11348 10810 11376 11698
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11624 10742 11652 13806
rect 11716 12918 11744 18294
rect 11900 17678 11928 19314
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 11992 18970 12020 19246
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11992 18426 12020 18906
rect 12084 18630 12112 19110
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 12084 17678 12112 18566
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 12084 16794 12112 17614
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11808 15706 11836 16186
rect 12084 15978 12112 16730
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 12072 15972 12124 15978
rect 12072 15914 12124 15920
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11808 12986 11836 15642
rect 11900 15609 11928 15914
rect 11886 15600 11942 15609
rect 11886 15535 11942 15544
rect 12176 15502 12204 19343
rect 12268 17882 12296 20266
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12544 20058 12572 20198
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 13096 19854 13124 20742
rect 13464 20058 13492 21490
rect 13556 21486 13584 22510
rect 13648 21894 13676 22578
rect 14175 22332 14483 22341
rect 14175 22330 14181 22332
rect 14237 22330 14261 22332
rect 14317 22330 14341 22332
rect 14397 22330 14421 22332
rect 14477 22330 14483 22332
rect 14237 22278 14239 22330
rect 14419 22278 14421 22330
rect 14175 22276 14181 22278
rect 14237 22276 14261 22278
rect 14317 22276 14341 22278
rect 14397 22276 14421 22278
rect 14477 22276 14483 22278
rect 14175 22267 14483 22276
rect 14280 21956 14332 21962
rect 14280 21898 14332 21904
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13648 21554 13676 21830
rect 13740 21690 13768 21830
rect 14292 21690 14320 21898
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 14835 21788 15143 21797
rect 14835 21786 14841 21788
rect 14897 21786 14921 21788
rect 14977 21786 15001 21788
rect 15057 21786 15081 21788
rect 15137 21786 15143 21788
rect 14897 21734 14899 21786
rect 15079 21734 15081 21786
rect 14835 21732 14841 21734
rect 14897 21732 14921 21734
rect 14977 21732 15001 21734
rect 15057 21732 15081 21734
rect 15137 21732 15143 21734
rect 14835 21723 15143 21732
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 15304 21622 15332 21830
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 15292 21616 15344 21622
rect 15292 21558 15344 21564
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 13556 21146 13584 21422
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 12912 19514 12940 19790
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12636 18698 12664 19314
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12452 18222 12480 18634
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12256 17128 12308 17134
rect 12452 17116 12480 17478
rect 12544 17338 12572 18226
rect 12636 17678 12664 18294
rect 12820 18222 12848 18566
rect 13004 18290 13032 19382
rect 13188 18426 13216 19790
rect 13280 19514 13308 19790
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13372 19446 13400 19858
rect 13360 19440 13412 19446
rect 13360 19382 13412 19388
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13556 18630 13584 19314
rect 14016 18952 14044 21422
rect 14108 21146 14136 21422
rect 15016 21412 15068 21418
rect 15016 21354 15068 21360
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14175 21244 14483 21253
rect 14175 21242 14181 21244
rect 14237 21242 14261 21244
rect 14317 21242 14341 21244
rect 14397 21242 14421 21244
rect 14477 21242 14483 21244
rect 14237 21190 14239 21242
rect 14419 21190 14421 21242
rect 14175 21188 14181 21190
rect 14237 21188 14261 21190
rect 14317 21188 14341 21190
rect 14397 21188 14421 21190
rect 14477 21188 14483 21190
rect 14175 21179 14483 21188
rect 14936 21146 14964 21286
rect 15028 21146 15056 21354
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 14835 20700 15143 20709
rect 14835 20698 14841 20700
rect 14897 20698 14921 20700
rect 14977 20698 15001 20700
rect 15057 20698 15081 20700
rect 15137 20698 15143 20700
rect 14897 20646 14899 20698
rect 15079 20646 15081 20698
rect 14835 20644 14841 20646
rect 14897 20644 14921 20646
rect 14977 20644 15001 20646
rect 15057 20644 15081 20646
rect 15137 20644 15143 20646
rect 14835 20635 15143 20644
rect 15212 20466 15240 21422
rect 15304 20602 15332 21422
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15488 21146 15516 21286
rect 15856 21146 15884 21490
rect 15476 21140 15528 21146
rect 15476 21082 15528 21088
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 16040 21078 16068 21490
rect 16132 21146 16160 21490
rect 16304 21344 16356 21350
rect 16302 21312 16304 21321
rect 16356 21312 16358 21321
rect 16302 21247 16358 21256
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 15568 21072 15620 21078
rect 15568 21014 15620 21020
rect 16028 21072 16080 21078
rect 16028 21014 16080 21020
rect 15580 20942 15608 21014
rect 15752 21004 15804 21010
rect 15752 20946 15804 20952
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 14175 20156 14483 20165
rect 14175 20154 14181 20156
rect 14237 20154 14261 20156
rect 14317 20154 14341 20156
rect 14397 20154 14421 20156
rect 14477 20154 14483 20156
rect 14237 20102 14239 20154
rect 14419 20102 14421 20154
rect 14175 20100 14181 20102
rect 14237 20100 14261 20102
rect 14317 20100 14341 20102
rect 14397 20100 14421 20102
rect 14477 20100 14483 20102
rect 14175 20091 14483 20100
rect 15212 19854 15240 20402
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15396 19786 15424 20402
rect 15488 20262 15516 20742
rect 15580 20602 15608 20878
rect 15764 20806 15792 20946
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 16408 20466 16436 21082
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15764 20058 15792 20402
rect 16132 20346 16160 20402
rect 16040 20318 16160 20346
rect 16212 20392 16264 20398
rect 16212 20334 16264 20340
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 14835 19612 15143 19621
rect 14835 19610 14841 19612
rect 14897 19610 14921 19612
rect 14977 19610 15001 19612
rect 15057 19610 15081 19612
rect 15137 19610 15143 19612
rect 14897 19558 14899 19610
rect 15079 19558 15081 19610
rect 14835 19556 14841 19558
rect 14897 19556 14921 19558
rect 14977 19556 15001 19558
rect 15057 19556 15081 19558
rect 15137 19556 15143 19558
rect 14835 19547 15143 19556
rect 14175 19068 14483 19077
rect 14175 19066 14181 19068
rect 14237 19066 14261 19068
rect 14317 19066 14341 19068
rect 14397 19066 14421 19068
rect 14477 19066 14483 19068
rect 14237 19014 14239 19066
rect 14419 19014 14421 19066
rect 14175 19012 14181 19014
rect 14237 19012 14261 19014
rect 14317 19012 14341 19014
rect 14397 19012 14421 19014
rect 14477 19012 14483 19014
rect 14175 19003 14483 19012
rect 13924 18924 14044 18952
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13556 18290 13584 18566
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 13740 17814 13768 18226
rect 13728 17808 13780 17814
rect 13728 17750 13780 17756
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13268 17604 13320 17610
rect 13268 17546 13320 17552
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 13004 17202 13032 17478
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12532 17128 12584 17134
rect 12452 17088 12532 17116
rect 12256 17070 12308 17076
rect 12532 17070 12584 17076
rect 12268 15910 12296 17070
rect 12820 16794 12848 17138
rect 12912 16794 12940 17138
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 12624 16720 12676 16726
rect 12624 16662 12676 16668
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12360 15570 12388 16390
rect 12452 15978 12480 16594
rect 12636 16182 12664 16662
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 12728 16114 12756 16526
rect 13004 16522 13032 16934
rect 13280 16658 13308 17546
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 12992 16516 13044 16522
rect 12992 16458 13044 16464
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12820 16114 12848 16390
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12900 15700 12952 15706
rect 12952 15660 13032 15688
rect 12900 15642 12952 15648
rect 13004 15570 13032 15660
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12176 14414 12204 15438
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 12820 15162 12848 15302
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 13096 14414 13124 15302
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11900 12102 11928 14350
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 14074 12664 14214
rect 13188 14074 13216 16526
rect 13280 16046 13308 16594
rect 13372 16522 13400 16934
rect 13464 16590 13492 17614
rect 13924 17270 13952 18924
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14004 18216 14056 18222
rect 14002 18184 14004 18193
rect 14056 18184 14058 18193
rect 14002 18119 14058 18128
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13360 16516 13412 16522
rect 13360 16458 13412 16464
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 13832 15162 13860 15574
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13740 14074 13768 14418
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12084 13394 12112 13806
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 11992 12442 12020 13194
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 13832 12306 13860 13126
rect 13924 12434 13952 17206
rect 14108 16046 14136 18702
rect 14372 18692 14424 18698
rect 14372 18634 14424 18640
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 14384 18426 14412 18634
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14568 18086 14596 18634
rect 14835 18524 15143 18533
rect 14835 18522 14841 18524
rect 14897 18522 14921 18524
rect 14977 18522 15001 18524
rect 15057 18522 15081 18524
rect 15137 18522 15143 18524
rect 14897 18470 14899 18522
rect 15079 18470 15081 18522
rect 14835 18468 14841 18470
rect 14897 18468 14921 18470
rect 14977 18468 15001 18470
rect 15057 18468 15081 18470
rect 15137 18468 15143 18470
rect 14835 18459 15143 18468
rect 15212 18358 15240 18634
rect 14740 18352 14792 18358
rect 14924 18352 14976 18358
rect 14792 18312 14872 18340
rect 14740 18294 14792 18300
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14660 18154 14688 18226
rect 14844 18222 14872 18312
rect 14924 18294 14976 18300
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14648 18148 14700 18154
rect 14648 18090 14700 18096
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14175 17980 14483 17989
rect 14175 17978 14181 17980
rect 14237 17978 14261 17980
rect 14317 17978 14341 17980
rect 14397 17978 14421 17980
rect 14477 17978 14483 17980
rect 14237 17926 14239 17978
rect 14419 17926 14421 17978
rect 14175 17924 14181 17926
rect 14237 17924 14261 17926
rect 14317 17924 14341 17926
rect 14397 17924 14421 17926
rect 14477 17924 14483 17926
rect 14175 17915 14483 17924
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14568 17270 14596 17546
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14660 17338 14688 17478
rect 14752 17338 14780 18022
rect 14844 17746 14872 18158
rect 14936 18086 14964 18294
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 14835 17436 15143 17445
rect 14835 17434 14841 17436
rect 14897 17434 14921 17436
rect 14977 17434 15001 17436
rect 15057 17434 15081 17436
rect 15137 17434 15143 17436
rect 14897 17382 14899 17434
rect 15079 17382 15081 17434
rect 14835 17380 14841 17382
rect 14897 17380 14921 17382
rect 14977 17380 15001 17382
rect 15057 17380 15081 17382
rect 15137 17380 15143 17382
rect 14835 17371 15143 17380
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 14175 16892 14483 16901
rect 14175 16890 14181 16892
rect 14237 16890 14261 16892
rect 14317 16890 14341 16892
rect 14397 16890 14421 16892
rect 14477 16890 14483 16892
rect 14237 16838 14239 16890
rect 14419 16838 14421 16890
rect 14175 16836 14181 16838
rect 14237 16836 14261 16838
rect 14317 16836 14341 16838
rect 14397 16836 14421 16838
rect 14477 16836 14483 16838
rect 14175 16827 14483 16836
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14476 16114 14504 16390
rect 14568 16266 14596 17206
rect 14660 16794 14688 17274
rect 15304 17202 15332 17614
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14568 16238 14688 16266
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14108 15094 14136 15982
rect 14175 15804 14483 15813
rect 14175 15802 14181 15804
rect 14237 15802 14261 15804
rect 14317 15802 14341 15804
rect 14397 15802 14421 15804
rect 14477 15802 14483 15804
rect 14237 15750 14239 15802
rect 14419 15750 14421 15802
rect 14175 15748 14181 15750
rect 14237 15748 14261 15750
rect 14317 15748 14341 15750
rect 14397 15748 14421 15750
rect 14477 15748 14483 15750
rect 14175 15739 14483 15748
rect 14568 15706 14596 16118
rect 14660 16114 14688 16238
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14292 15162 14320 15438
rect 14660 15314 14688 16050
rect 14752 15722 14780 16390
rect 14835 16348 15143 16357
rect 14835 16346 14841 16348
rect 14897 16346 14921 16348
rect 14977 16346 15001 16348
rect 15057 16346 15081 16348
rect 15137 16346 15143 16348
rect 14897 16294 14899 16346
rect 15079 16294 15081 16346
rect 14835 16292 14841 16294
rect 14897 16292 14921 16294
rect 14977 16292 15001 16294
rect 15057 16292 15081 16294
rect 15137 16292 15143 16294
rect 14835 16283 15143 16292
rect 15212 16250 15240 17002
rect 15304 16794 15332 17138
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 14924 16108 14976 16114
rect 14844 16068 14924 16096
rect 14844 15910 14872 16068
rect 14924 16050 14976 16056
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14752 15694 14964 15722
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14844 15348 14872 15438
rect 14936 15434 14964 15694
rect 15212 15502 15240 16186
rect 15290 15600 15346 15609
rect 15290 15535 15346 15544
rect 15304 15502 15332 15535
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 14752 15320 14872 15348
rect 14752 15314 14780 15320
rect 14660 15286 14780 15314
rect 14660 15162 14688 15286
rect 14835 15260 15143 15269
rect 14835 15258 14841 15260
rect 14897 15258 14921 15260
rect 14977 15258 15001 15260
rect 15057 15258 15081 15260
rect 15137 15258 15143 15260
rect 14897 15206 14899 15258
rect 15079 15206 15081 15258
rect 14835 15204 14841 15206
rect 14897 15204 14921 15206
rect 14977 15204 15001 15206
rect 15057 15204 15081 15206
rect 15137 15204 15143 15206
rect 14835 15195 15143 15204
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14175 14716 14483 14725
rect 14175 14714 14181 14716
rect 14237 14714 14261 14716
rect 14317 14714 14341 14716
rect 14397 14714 14421 14716
rect 14477 14714 14483 14716
rect 14237 14662 14239 14714
rect 14419 14662 14421 14714
rect 14175 14660 14181 14662
rect 14237 14660 14261 14662
rect 14317 14660 14341 14662
rect 14397 14660 14421 14662
rect 14477 14660 14483 14662
rect 14175 14651 14483 14660
rect 14568 14618 14596 14758
rect 15212 14618 15240 14962
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14384 14074 14412 14214
rect 14476 14074 14504 14214
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14568 13734 14596 14554
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14660 13802 14688 14350
rect 14835 14172 15143 14181
rect 14835 14170 14841 14172
rect 14897 14170 14921 14172
rect 14977 14170 15001 14172
rect 15057 14170 15081 14172
rect 15137 14170 15143 14172
rect 14897 14118 14899 14170
rect 15079 14118 15081 14170
rect 14835 14116 14841 14118
rect 14897 14116 14921 14118
rect 14977 14116 15001 14118
rect 15057 14116 15081 14118
rect 15137 14116 15143 14118
rect 14835 14107 15143 14116
rect 15212 14074 15240 14554
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 15304 14074 15332 14418
rect 15396 14074 15424 19722
rect 16040 19718 16068 20318
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16132 19938 16160 20198
rect 16224 20058 16252 20334
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16408 20058 16436 20198
rect 16212 20052 16264 20058
rect 16212 19994 16264 20000
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16132 19910 16252 19938
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15580 18193 15608 18770
rect 15566 18184 15622 18193
rect 15566 18119 15622 18128
rect 15580 17542 15608 18119
rect 16040 17882 16068 19654
rect 16224 19174 16252 19910
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16316 19514 16344 19790
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16316 19378 16344 19450
rect 16592 19417 16620 21626
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16684 20330 16712 21490
rect 16776 21434 16804 22578
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 16960 21962 16988 22374
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16776 21406 16896 21434
rect 16868 21350 16896 21406
rect 16948 21412 17000 21418
rect 16948 21354 17000 21360
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16856 21344 16908 21350
rect 16960 21321 16988 21354
rect 16856 21286 16908 21292
rect 16946 21312 17002 21321
rect 16776 21146 16804 21286
rect 16946 21247 17002 21256
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16672 20324 16724 20330
rect 16672 20266 16724 20272
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16578 19408 16634 19417
rect 16304 19372 16356 19378
rect 16776 19378 16804 19654
rect 16578 19343 16634 19352
rect 16764 19372 16816 19378
rect 16304 19314 16356 19320
rect 16764 19314 16816 19320
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 16224 17678 16252 19110
rect 16316 18970 16344 19314
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16592 18902 16620 19246
rect 16960 18970 16988 20402
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17420 19378 17448 19994
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17604 19514 17632 19790
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 17052 19174 17080 19246
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17144 18970 17172 19110
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17144 18222 17172 18634
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17052 18086 17080 18158
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 16592 17678 16620 18022
rect 17052 17882 17080 18022
rect 17420 17882 17448 19314
rect 17776 18964 17828 18970
rect 17828 18924 18092 18952
rect 17776 18906 17828 18912
rect 18064 18834 18092 18924
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 18156 18766 18184 19654
rect 19076 19378 19104 21966
rect 19352 19938 19380 22374
rect 19465 22332 19773 22341
rect 19465 22330 19471 22332
rect 19527 22330 19551 22332
rect 19607 22330 19631 22332
rect 19687 22330 19711 22332
rect 19767 22330 19773 22332
rect 19527 22278 19529 22330
rect 19709 22278 19711 22330
rect 19465 22276 19471 22278
rect 19527 22276 19551 22278
rect 19607 22276 19631 22278
rect 19687 22276 19711 22278
rect 19767 22276 19773 22278
rect 19465 22267 19773 22276
rect 20125 21788 20433 21797
rect 20125 21786 20131 21788
rect 20187 21786 20211 21788
rect 20267 21786 20291 21788
rect 20347 21786 20371 21788
rect 20427 21786 20433 21788
rect 20187 21734 20189 21786
rect 20369 21734 20371 21786
rect 20125 21732 20131 21734
rect 20187 21732 20211 21734
rect 20267 21732 20291 21734
rect 20347 21732 20371 21734
rect 20427 21732 20433 21734
rect 20125 21723 20433 21732
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 19465 21244 19773 21253
rect 19465 21242 19471 21244
rect 19527 21242 19551 21244
rect 19607 21242 19631 21244
rect 19687 21242 19711 21244
rect 19767 21242 19773 21244
rect 19527 21190 19529 21242
rect 19709 21190 19711 21242
rect 19465 21188 19471 21190
rect 19527 21188 19551 21190
rect 19607 21188 19631 21190
rect 19687 21188 19711 21190
rect 19767 21188 19773 21190
rect 19465 21179 19773 21188
rect 20125 20700 20433 20709
rect 20125 20698 20131 20700
rect 20187 20698 20211 20700
rect 20267 20698 20291 20700
rect 20347 20698 20371 20700
rect 20427 20698 20433 20700
rect 20187 20646 20189 20698
rect 20369 20646 20371 20698
rect 20125 20644 20131 20646
rect 20187 20644 20211 20646
rect 20267 20644 20291 20646
rect 20347 20644 20371 20646
rect 20427 20644 20433 20646
rect 20125 20635 20433 20644
rect 20640 20602 20668 21286
rect 22204 21185 22232 21490
rect 22190 21176 22246 21185
rect 22190 21111 22246 21120
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 19465 20156 19773 20165
rect 19465 20154 19471 20156
rect 19527 20154 19551 20156
rect 19607 20154 19631 20156
rect 19687 20154 19711 20156
rect 19767 20154 19773 20156
rect 19527 20102 19529 20154
rect 19709 20102 19711 20154
rect 19465 20100 19471 20102
rect 19527 20100 19551 20102
rect 19607 20100 19631 20102
rect 19687 20100 19711 20102
rect 19767 20100 19773 20102
rect 19465 20091 19773 20100
rect 20180 19990 20208 20198
rect 20548 20058 20576 20198
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20168 19984 20220 19990
rect 19352 19910 19472 19938
rect 20168 19926 20220 19932
rect 19444 19854 19472 19910
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 19260 19514 19288 19654
rect 20125 19612 20433 19621
rect 20125 19610 20131 19612
rect 20187 19610 20211 19612
rect 20267 19610 20291 19612
rect 20347 19610 20371 19612
rect 20427 19610 20433 19612
rect 20187 19558 20189 19610
rect 20369 19558 20371 19610
rect 20125 19556 20131 19558
rect 20187 19556 20211 19558
rect 20267 19556 20291 19558
rect 20347 19556 20371 19558
rect 20427 19556 20433 19558
rect 20125 19547 20433 19556
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18340 18970 18368 19314
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 19352 18766 19380 19246
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19465 19068 19773 19077
rect 19465 19066 19471 19068
rect 19527 19066 19551 19068
rect 19607 19066 19631 19068
rect 19687 19066 19711 19068
rect 19767 19066 19773 19068
rect 19527 19014 19529 19066
rect 19709 19014 19711 19066
rect 19465 19012 19471 19014
rect 19527 19012 19551 19014
rect 19607 19012 19631 19014
rect 19687 19012 19711 19014
rect 19767 19012 19773 19014
rect 19465 19003 19773 19012
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17512 18358 17540 18634
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15580 17270 15608 17478
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15488 16658 15516 17138
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15488 16250 15516 16594
rect 15580 16590 15608 17206
rect 16224 17202 16252 17614
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16960 17134 16988 17614
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15580 15162 15608 16526
rect 16960 16114 16988 17070
rect 18524 16794 18552 17138
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 19260 16658 19288 18566
rect 19352 17270 19380 18702
rect 19904 18698 19932 19110
rect 19892 18692 19944 18698
rect 19892 18634 19944 18640
rect 20125 18524 20433 18533
rect 20125 18522 20131 18524
rect 20187 18522 20211 18524
rect 20267 18522 20291 18524
rect 20347 18522 20371 18524
rect 20427 18522 20433 18524
rect 20187 18470 20189 18522
rect 20369 18470 20371 18522
rect 20125 18468 20131 18470
rect 20187 18468 20211 18470
rect 20267 18468 20291 18470
rect 20347 18468 20371 18470
rect 20427 18468 20433 18470
rect 20125 18459 20433 18468
rect 19465 17980 19773 17989
rect 19465 17978 19471 17980
rect 19527 17978 19551 17980
rect 19607 17978 19631 17980
rect 19687 17978 19711 17980
rect 19767 17978 19773 17980
rect 19527 17926 19529 17978
rect 19709 17926 19711 17978
rect 19465 17924 19471 17926
rect 19527 17924 19551 17926
rect 19607 17924 19631 17926
rect 19687 17924 19711 17926
rect 19767 17924 19773 17926
rect 19465 17915 19773 17924
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19465 16892 19773 16901
rect 19465 16890 19471 16892
rect 19527 16890 19551 16892
rect 19607 16890 19631 16892
rect 19687 16890 19711 16892
rect 19767 16890 19773 16892
rect 19527 16838 19529 16890
rect 19709 16838 19711 16890
rect 19465 16836 19471 16838
rect 19527 16836 19551 16838
rect 19607 16836 19631 16838
rect 19687 16836 19711 16838
rect 19767 16836 19773 16838
rect 19465 16827 19773 16836
rect 19812 16794 19840 17614
rect 19892 17536 19944 17542
rect 19892 17478 19944 17484
rect 19904 17338 19932 17478
rect 20125 17436 20433 17445
rect 20125 17434 20131 17436
rect 20187 17434 20211 17436
rect 20267 17434 20291 17436
rect 20347 17434 20371 17436
rect 20427 17434 20433 17436
rect 20187 17382 20189 17434
rect 20369 17382 20371 17434
rect 20125 17380 20131 17382
rect 20187 17380 20211 17382
rect 20267 17380 20291 17382
rect 20347 17380 20371 17382
rect 20427 17380 20433 17382
rect 20125 17371 20433 17380
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17236 16114 17264 16390
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 16960 15706 16988 16050
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14175 13628 14483 13637
rect 14175 13626 14181 13628
rect 14237 13626 14261 13628
rect 14317 13626 14341 13628
rect 14397 13626 14421 13628
rect 14477 13626 14483 13628
rect 14237 13574 14239 13626
rect 14419 13574 14421 13626
rect 14175 13572 14181 13574
rect 14237 13572 14261 13574
rect 14317 13572 14341 13574
rect 14397 13572 14421 13574
rect 14477 13572 14483 13574
rect 14175 13563 14483 13572
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14568 12918 14596 13126
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14660 12714 14688 13738
rect 14835 13084 15143 13093
rect 14835 13082 14841 13084
rect 14897 13082 14921 13084
rect 14977 13082 15001 13084
rect 15057 13082 15081 13084
rect 15137 13082 15143 13084
rect 14897 13030 14899 13082
rect 15079 13030 15081 13082
rect 14835 13028 14841 13030
rect 14897 13028 14921 13030
rect 14977 13028 15001 13030
rect 15057 13028 15081 13030
rect 15137 13028 15143 13030
rect 14835 13019 15143 13028
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14175 12540 14483 12549
rect 14175 12538 14181 12540
rect 14237 12538 14261 12540
rect 14317 12538 14341 12540
rect 14397 12538 14421 12540
rect 14477 12538 14483 12540
rect 14237 12486 14239 12538
rect 14419 12486 14421 12538
rect 14175 12484 14181 12486
rect 14237 12484 14261 12486
rect 14317 12484 14341 12486
rect 14397 12484 14421 12486
rect 14477 12484 14483 12486
rect 14175 12475 14483 12484
rect 13924 12406 14412 12434
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13924 12102 13952 12406
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13004 11898 13032 12038
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 14016 11830 14044 12038
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11624 10062 11652 10678
rect 11808 10674 11836 11494
rect 12268 11014 12296 11630
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12360 11082 12388 11494
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 12268 10538 12296 10950
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 12084 10266 12112 10406
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 12268 9994 12296 10474
rect 12544 10266 12572 11698
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12636 10674 12664 11290
rect 12820 10810 12848 11562
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12636 10062 12664 10610
rect 12912 10266 12940 11698
rect 14384 11694 14412 12406
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14372 11688 14424 11694
rect 14372 11630 14424 11636
rect 14175 11452 14483 11461
rect 14175 11450 14181 11452
rect 14237 11450 14261 11452
rect 14317 11450 14341 11452
rect 14397 11450 14421 11452
rect 14477 11450 14483 11452
rect 14237 11398 14239 11450
rect 14419 11398 14421 11450
rect 14175 11396 14181 11398
rect 14237 11396 14261 11398
rect 14317 11396 14341 11398
rect 14397 11396 14421 11398
rect 14477 11396 14483 11398
rect 14175 11387 14483 11396
rect 14568 11354 14596 12174
rect 14648 11824 14700 11830
rect 14648 11766 14700 11772
rect 14660 11354 14688 11766
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13556 11014 13584 11154
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12624 10056 12676 10062
rect 13464 10044 13492 10542
rect 13556 10248 13584 10950
rect 13648 10606 13676 10950
rect 13832 10674 13860 10950
rect 14568 10810 14596 11018
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 14175 10364 14483 10373
rect 14175 10362 14181 10364
rect 14237 10362 14261 10364
rect 14317 10362 14341 10364
rect 14397 10362 14421 10364
rect 14477 10362 14483 10364
rect 14237 10310 14239 10362
rect 14419 10310 14421 10362
rect 14175 10308 14181 10310
rect 14237 10308 14261 10310
rect 14317 10308 14341 10310
rect 14397 10308 14421 10310
rect 14477 10308 14483 10310
rect 14175 10299 14483 10308
rect 13636 10260 13688 10266
rect 13556 10220 13636 10248
rect 13636 10202 13688 10208
rect 13544 10056 13596 10062
rect 13464 10016 13544 10044
rect 12624 9998 12676 10004
rect 13544 9998 13596 10004
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12360 9722 12388 9998
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11428 9172 11480 9178
rect 11256 9132 11428 9160
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11164 8922 11192 9046
rect 11256 9042 11284 9132
rect 11428 9114 11480 9120
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11348 8922 11376 8978
rect 11164 8894 11376 8922
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8362 11100 8774
rect 11336 8628 11388 8634
rect 11440 8616 11468 8978
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11388 8588 11468 8616
rect 11336 8570 11388 8576
rect 11532 8537 11560 8910
rect 11518 8528 11574 8537
rect 11624 8498 11652 9318
rect 11808 9178 11836 9522
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11900 9178 11928 9454
rect 13556 9178 13584 9998
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9586 14136 9862
rect 14384 9654 14412 9998
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14175 9276 14483 9285
rect 14175 9274 14181 9276
rect 14237 9274 14261 9276
rect 14317 9274 14341 9276
rect 14397 9274 14421 9276
rect 14477 9274 14483 9276
rect 14237 9222 14239 9274
rect 14419 9222 14421 9274
rect 14175 9220 14181 9222
rect 14237 9220 14261 9222
rect 14317 9220 14341 9222
rect 14397 9220 14421 9222
rect 14477 9220 14483 9222
rect 14175 9211 14483 9220
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 11716 8634 11744 8910
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11518 8463 11574 8472
rect 11612 8492 11664 8498
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10888 8078 11100 8106
rect 11440 8090 11468 8366
rect 11072 7970 11100 8078
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11072 7942 11192 7970
rect 11164 6866 11192 7942
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11164 6202 11192 6802
rect 11532 6458 11560 8463
rect 11612 8434 11664 8440
rect 11716 7546 11744 8570
rect 12084 8090 12112 8910
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12360 7886 12388 8774
rect 12728 8634 12756 8910
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 13464 8362 13492 8774
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13648 8090 13676 8434
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11992 7546 12020 7754
rect 12452 7546 12480 7822
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 12084 6798 12112 7278
rect 12544 7002 12572 7822
rect 12636 7206 12664 7822
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11900 6458 11928 6734
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 12084 6322 12112 6734
rect 12636 6390 12664 7142
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 11164 6174 11284 6202
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10612 5370 10640 5714
rect 11164 5710 11192 6054
rect 11152 5704 11204 5710
rect 11150 5672 11152 5681
rect 11204 5672 11206 5681
rect 11150 5607 11206 5616
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10704 3670 10732 3878
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10600 3528 10652 3534
rect 10876 3528 10928 3534
rect 10600 3470 10652 3476
rect 10796 3476 10876 3482
rect 10796 3470 10928 3476
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 9416 3176 9444 3334
rect 9545 3292 9853 3301
rect 9545 3290 9551 3292
rect 9607 3290 9631 3292
rect 9687 3290 9711 3292
rect 9767 3290 9791 3292
rect 9847 3290 9853 3292
rect 9607 3238 9609 3290
rect 9789 3238 9791 3290
rect 9545 3236 9551 3238
rect 9607 3236 9631 3238
rect 9687 3236 9711 3238
rect 9767 3236 9791 3238
rect 9847 3236 9853 3238
rect 9545 3227 9853 3236
rect 10060 3194 10088 3334
rect 10048 3188 10100 3194
rect 9416 3148 9536 3176
rect 9508 3058 9536 3148
rect 10048 3130 10100 3136
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 10612 2922 10640 3470
rect 10796 3454 10916 3470
rect 10796 3126 10824 3454
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 10888 2922 10916 3334
rect 11072 3058 11100 3878
rect 11256 3738 11284 6174
rect 12084 5710 12112 6258
rect 13280 6186 13308 6326
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 13268 6180 13320 6186
rect 13268 6122 13320 6128
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12176 5642 12204 6122
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 13096 5914 13124 6054
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13740 5710 13768 8230
rect 13832 8022 13860 8230
rect 14108 8090 14136 8434
rect 14175 8188 14483 8197
rect 14175 8186 14181 8188
rect 14237 8186 14261 8188
rect 14317 8186 14341 8188
rect 14397 8186 14421 8188
rect 14477 8186 14483 8188
rect 14237 8134 14239 8186
rect 14419 8134 14421 8186
rect 14175 8132 14181 8134
rect 14237 8132 14261 8134
rect 14317 8132 14341 8134
rect 14397 8132 14421 8134
rect 14477 8132 14483 8134
rect 14175 8123 14483 8132
rect 14568 8090 14596 9590
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14568 7478 14596 7686
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13924 6866 13952 7346
rect 14175 7100 14483 7109
rect 14175 7098 14181 7100
rect 14237 7098 14261 7100
rect 14317 7098 14341 7100
rect 14397 7098 14421 7100
rect 14477 7098 14483 7100
rect 14237 7046 14239 7098
rect 14419 7046 14421 7098
rect 14175 7044 14181 7046
rect 14237 7044 14261 7046
rect 14317 7044 14341 7046
rect 14397 7044 14421 7046
rect 14477 7044 14483 7046
rect 14175 7035 14483 7044
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13924 6458 13952 6802
rect 14568 6798 14596 7414
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14660 6662 14688 7346
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14108 6458 14136 6598
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14175 6012 14483 6021
rect 14175 6010 14181 6012
rect 14237 6010 14261 6012
rect 14317 6010 14341 6012
rect 14397 6010 14421 6012
rect 14477 6010 14483 6012
rect 14237 5958 14239 6010
rect 14419 5958 14421 6010
rect 14175 5956 14181 5958
rect 14237 5956 14261 5958
rect 14317 5956 14341 5958
rect 14397 5956 14421 5958
rect 14477 5956 14483 5958
rect 14175 5947 14483 5956
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 13280 5030 13308 5646
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11716 4282 11744 4694
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11716 4010 11744 4082
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11164 3194 11192 3470
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11256 3058 11284 3674
rect 11808 3126 11836 3878
rect 12636 3738 12664 4150
rect 12912 3942 12940 4966
rect 13832 4826 13860 5578
rect 14660 5370 14688 6598
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14752 5302 14780 12854
rect 15304 12850 15332 13874
rect 15488 13734 15516 14350
rect 15580 14074 15608 14962
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13530 15516 13670
rect 15580 13530 15608 13806
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 13530 15700 13670
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15396 12782 15424 13126
rect 15672 12850 15700 13466
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 14835 11996 15143 12005
rect 14835 11994 14841 11996
rect 14897 11994 14921 11996
rect 14977 11994 15001 11996
rect 15057 11994 15081 11996
rect 15137 11994 15143 11996
rect 14897 11942 14899 11994
rect 15079 11942 15081 11994
rect 14835 11940 14841 11942
rect 14897 11940 14921 11942
rect 14977 11940 15001 11942
rect 15057 11940 15081 11942
rect 15137 11940 15143 11942
rect 14835 11931 15143 11940
rect 15764 11898 15792 15370
rect 16684 15162 16712 15438
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 16960 15026 16988 15642
rect 17604 15434 17632 16526
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16304 14544 16356 14550
rect 16304 14486 16356 14492
rect 16316 14074 16344 14486
rect 16960 14482 16988 14962
rect 18064 14618 18092 16390
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18248 14958 18276 15438
rect 18340 15366 18368 16594
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 19076 16250 19104 16526
rect 19708 16448 19760 16454
rect 19708 16390 19760 16396
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19614 16008 19670 16017
rect 19614 15943 19616 15952
rect 19668 15943 19670 15952
rect 19616 15914 19668 15920
rect 19720 15910 19748 16390
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 18420 15904 18472 15910
rect 19432 15904 19484 15910
rect 18420 15846 18472 15852
rect 19352 15864 19432 15892
rect 18432 15502 18460 15846
rect 19352 15688 19380 15864
rect 19432 15846 19484 15852
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 19465 15804 19773 15813
rect 19465 15802 19471 15804
rect 19527 15802 19551 15804
rect 19607 15802 19631 15804
rect 19687 15802 19711 15804
rect 19767 15802 19773 15804
rect 19527 15750 19529 15802
rect 19709 15750 19711 15802
rect 19465 15748 19471 15750
rect 19527 15748 19551 15750
rect 19607 15748 19631 15750
rect 19687 15748 19711 15750
rect 19767 15748 19773 15750
rect 19465 15739 19773 15748
rect 19432 15700 19484 15706
rect 19352 15660 19432 15688
rect 19432 15642 19484 15648
rect 19338 15600 19394 15609
rect 19338 15535 19394 15544
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18340 15026 18368 15302
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18432 14822 18460 15438
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18616 15094 18644 15302
rect 18892 15162 18920 15302
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18616 14618 18644 15030
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16776 13938 16804 14350
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 16960 14074 16988 14214
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16500 12986 16528 13194
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 16040 12434 16068 12786
rect 16040 12406 16160 12434
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15948 11830 15976 12106
rect 15936 11824 15988 11830
rect 15936 11766 15988 11772
rect 15292 11144 15344 11150
rect 15948 11098 15976 11766
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 15292 11086 15344 11092
rect 14835 10908 15143 10917
rect 14835 10906 14841 10908
rect 14897 10906 14921 10908
rect 14977 10906 15001 10908
rect 15057 10906 15081 10908
rect 15137 10906 15143 10908
rect 14897 10854 14899 10906
rect 15079 10854 15081 10906
rect 14835 10852 14841 10854
rect 14897 10852 14921 10854
rect 14977 10852 15001 10854
rect 15057 10852 15081 10854
rect 15137 10852 15143 10854
rect 14835 10843 15143 10852
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14844 10266 14872 10610
rect 15304 10470 15332 11086
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15856 11070 15976 11098
rect 15396 10674 15424 11018
rect 15672 10742 15700 11018
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 10266 15792 10406
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 14835 9820 15143 9829
rect 14835 9818 14841 9820
rect 14897 9818 14921 9820
rect 14977 9818 15001 9820
rect 15057 9818 15081 9820
rect 15137 9818 15143 9820
rect 14897 9766 14899 9818
rect 15079 9766 15081 9818
rect 14835 9764 14841 9766
rect 14897 9764 14921 9766
rect 14977 9764 15001 9766
rect 15057 9764 15081 9766
rect 15137 9764 15143 9766
rect 14835 9755 15143 9764
rect 15396 8974 15424 9998
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 14835 8732 15143 8741
rect 14835 8730 14841 8732
rect 14897 8730 14921 8732
rect 14977 8730 15001 8732
rect 15057 8730 15081 8732
rect 15137 8730 15143 8732
rect 14897 8678 14899 8730
rect 15079 8678 15081 8730
rect 14835 8676 14841 8678
rect 14897 8676 14921 8678
rect 14977 8676 15001 8678
rect 15057 8676 15081 8678
rect 15137 8676 15143 8678
rect 14835 8667 15143 8676
rect 15212 8090 15240 8842
rect 15396 8566 15424 8910
rect 15384 8560 15436 8566
rect 15384 8502 15436 8508
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 14835 7644 15143 7653
rect 14835 7642 14841 7644
rect 14897 7642 14921 7644
rect 14977 7642 15001 7644
rect 15057 7642 15081 7644
rect 15137 7642 15143 7644
rect 14897 7590 14899 7642
rect 15079 7590 15081 7642
rect 14835 7588 14841 7590
rect 14897 7588 14921 7590
rect 14977 7588 15001 7590
rect 15057 7588 15081 7590
rect 15137 7588 15143 7590
rect 14835 7579 15143 7588
rect 15304 7342 15332 8230
rect 15396 7954 15424 8502
rect 15856 8498 15884 11070
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 10810 15976 10950
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 16040 10690 16068 11698
rect 15948 10674 16068 10690
rect 15936 10668 16068 10674
rect 15988 10662 16068 10668
rect 15936 10610 15988 10616
rect 16040 9722 16068 10662
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16132 8974 16160 12406
rect 16776 11830 16804 13874
rect 17604 13802 17632 14282
rect 18616 13938 18644 14554
rect 19076 14074 19104 15438
rect 19352 15094 19380 15535
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19444 15026 19472 15302
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19628 14890 19656 15370
rect 19720 15162 19748 15370
rect 19812 15162 19840 16186
rect 19904 16114 19932 17138
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20088 16658 20116 16934
rect 20076 16652 20128 16658
rect 20076 16594 20128 16600
rect 20088 16561 20116 16594
rect 20074 16552 20130 16561
rect 20074 16487 20130 16496
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19996 16250 20024 16390
rect 20125 16348 20433 16357
rect 20125 16346 20131 16348
rect 20187 16346 20211 16348
rect 20267 16346 20291 16348
rect 20347 16346 20371 16348
rect 20427 16346 20433 16348
rect 20187 16294 20189 16346
rect 20369 16294 20371 16346
rect 20125 16292 20131 16294
rect 20187 16292 20211 16294
rect 20267 16292 20291 16294
rect 20347 16292 20371 16294
rect 20427 16292 20433 16294
rect 20125 16283 20433 16292
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 19982 16144 20038 16153
rect 19892 16108 19944 16114
rect 19982 16079 20038 16088
rect 19892 16050 19944 16056
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19904 15638 19932 15846
rect 19996 15706 20024 16079
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20272 15706 20300 15846
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 19892 15632 19944 15638
rect 19892 15574 19944 15580
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19904 14958 19932 15438
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19616 14884 19668 14890
rect 19616 14826 19668 14832
rect 19260 14618 19288 14826
rect 19996 14822 20024 15642
rect 20364 15434 20392 16186
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20352 15428 20404 15434
rect 20352 15370 20404 15376
rect 20125 15260 20433 15269
rect 20125 15258 20131 15260
rect 20187 15258 20211 15260
rect 20267 15258 20291 15260
rect 20347 15258 20371 15260
rect 20427 15258 20433 15260
rect 20187 15206 20189 15258
rect 20369 15206 20371 15258
rect 20125 15204 20131 15206
rect 20187 15204 20211 15206
rect 20267 15204 20291 15206
rect 20347 15204 20371 15206
rect 20427 15204 20433 15206
rect 20125 15195 20433 15204
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19352 14618 19380 14758
rect 19465 14716 19773 14725
rect 19465 14714 19471 14716
rect 19527 14714 19551 14716
rect 19607 14714 19631 14716
rect 19687 14714 19711 14716
rect 19767 14714 19773 14716
rect 19527 14662 19529 14714
rect 19709 14662 19711 14714
rect 19465 14660 19471 14662
rect 19527 14660 19551 14662
rect 19607 14660 19631 14662
rect 19687 14660 19711 14662
rect 19767 14660 19773 14662
rect 19465 14651 19773 14660
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 19465 13628 19773 13637
rect 19465 13626 19471 13628
rect 19527 13626 19551 13628
rect 19607 13626 19631 13628
rect 19687 13626 19711 13628
rect 19767 13626 19773 13628
rect 19527 13574 19529 13626
rect 19709 13574 19711 13626
rect 19465 13572 19471 13574
rect 19527 13572 19551 13574
rect 19607 13572 19631 13574
rect 19687 13572 19711 13574
rect 19767 13572 19773 13574
rect 19465 13563 19773 13572
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17512 12434 17540 12582
rect 17604 12442 17632 13262
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 18064 12850 18092 13194
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17328 12406 17540 12434
rect 17592 12436 17644 12442
rect 17328 12238 17356 12406
rect 17592 12378 17644 12384
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 17604 11762 17632 12378
rect 18708 12374 18736 13262
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16500 10810 16528 11494
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16500 10198 16528 10542
rect 16488 10192 16540 10198
rect 16488 10134 16540 10140
rect 16684 9722 16712 10610
rect 16868 10470 16896 11018
rect 17236 11014 17264 11630
rect 17604 11218 17632 11698
rect 19168 11354 19196 12038
rect 19260 11830 19288 13126
rect 19720 12782 19748 13126
rect 19812 12918 19840 13126
rect 19800 12912 19852 12918
rect 19800 12854 19852 12860
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19465 12540 19773 12549
rect 19465 12538 19471 12540
rect 19527 12538 19551 12540
rect 19607 12538 19631 12540
rect 19687 12538 19711 12540
rect 19767 12538 19773 12540
rect 19527 12486 19529 12538
rect 19709 12486 19711 12538
rect 19465 12484 19471 12486
rect 19527 12484 19551 12486
rect 19607 12484 19631 12486
rect 19687 12484 19711 12486
rect 19767 12484 19773 12486
rect 19465 12475 19773 12484
rect 19904 12322 19932 14758
rect 20125 14172 20433 14181
rect 20125 14170 20131 14172
rect 20187 14170 20211 14172
rect 20267 14170 20291 14172
rect 20347 14170 20371 14172
rect 20427 14170 20433 14172
rect 20187 14118 20189 14170
rect 20369 14118 20371 14170
rect 20125 14116 20131 14118
rect 20187 14116 20211 14118
rect 20267 14116 20291 14118
rect 20347 14116 20371 14118
rect 20427 14116 20433 14118
rect 20125 14107 20433 14116
rect 20548 13938 20576 15438
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 19996 12986 20024 13874
rect 20272 13818 20300 13874
rect 20640 13818 20668 19654
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20916 16794 20944 17478
rect 21468 17338 21496 17614
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20732 15162 20760 16390
rect 21468 16250 21496 17274
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21652 16250 21680 16526
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21652 15502 21680 16186
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 20904 15428 20956 15434
rect 20904 15370 20956 15376
rect 20916 15162 20944 15370
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 20272 13790 20668 13818
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 13326 21404 13670
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 20125 13084 20433 13093
rect 20125 13082 20131 13084
rect 20187 13082 20211 13084
rect 20267 13082 20291 13084
rect 20347 13082 20371 13084
rect 20427 13082 20433 13084
rect 20187 13030 20189 13082
rect 20369 13030 20371 13082
rect 20125 13028 20131 13030
rect 20187 13028 20211 13030
rect 20267 13028 20291 13030
rect 20347 13028 20371 13030
rect 20427 13028 20433 13030
rect 20125 13019 20433 13028
rect 20640 12986 20668 13262
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 19996 12442 20024 12922
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19904 12294 20024 12322
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19248 11824 19300 11830
rect 19248 11766 19300 11772
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19260 11354 19288 11630
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19465 11452 19773 11461
rect 19465 11450 19471 11452
rect 19527 11450 19551 11452
rect 19607 11450 19631 11452
rect 19687 11450 19711 11452
rect 19767 11450 19773 11452
rect 19527 11398 19529 11450
rect 19709 11398 19711 11450
rect 19465 11396 19471 11398
rect 19527 11396 19551 11398
rect 19607 11396 19631 11398
rect 19687 11396 19711 11398
rect 19767 11396 19773 11398
rect 19465 11387 19773 11396
rect 19812 11354 19840 11494
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 18236 11212 18288 11218
rect 18236 11154 18288 11160
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17236 10810 17264 10950
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 18248 10674 18276 11154
rect 19352 10742 19380 11222
rect 19812 11014 19840 11290
rect 19904 11286 19932 12174
rect 19892 11280 19944 11286
rect 19892 11222 19944 11228
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 19465 10364 19773 10373
rect 19465 10362 19471 10364
rect 19527 10362 19551 10364
rect 19607 10362 19631 10364
rect 19687 10362 19711 10364
rect 19767 10362 19773 10364
rect 19527 10310 19529 10362
rect 19709 10310 19711 10362
rect 19465 10308 19471 10310
rect 19527 10308 19551 10310
rect 19607 10308 19631 10310
rect 19687 10308 19711 10310
rect 19767 10308 19773 10310
rect 19465 10299 19773 10308
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 17236 9518 17264 9862
rect 18432 9586 18460 9862
rect 19076 9722 19104 9998
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 16132 8634 16160 8910
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 15488 7886 15516 8230
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15856 6798 15884 8434
rect 16132 6866 16160 8570
rect 16592 8498 16620 8774
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 15844 6792 15896 6798
rect 15764 6740 15844 6746
rect 15764 6734 15896 6740
rect 15764 6718 15884 6734
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 14835 6556 15143 6565
rect 14835 6554 14841 6556
rect 14897 6554 14921 6556
rect 14977 6554 15001 6556
rect 15057 6554 15081 6556
rect 15137 6554 15143 6556
rect 14897 6502 14899 6554
rect 15079 6502 15081 6554
rect 14835 6500 14841 6502
rect 14897 6500 14921 6502
rect 14977 6500 15001 6502
rect 15057 6500 15081 6502
rect 15137 6500 15143 6502
rect 14835 6491 15143 6500
rect 15488 6458 15516 6598
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15304 5710 15332 6190
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15488 5914 15516 6054
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 14835 5468 15143 5477
rect 14835 5466 14841 5468
rect 14897 5466 14921 5468
rect 14977 5466 15001 5468
rect 15057 5466 15081 5468
rect 15137 5466 15143 5468
rect 14897 5414 14899 5466
rect 15079 5414 15081 5466
rect 14835 5412 14841 5414
rect 14897 5412 14921 5414
rect 14977 5412 15001 5414
rect 15057 5412 15081 5414
rect 15137 5412 15143 5414
rect 14835 5403 15143 5412
rect 14740 5296 14792 5302
rect 14740 5238 14792 5244
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 14175 4924 14483 4933
rect 14175 4922 14181 4924
rect 14237 4922 14261 4924
rect 14317 4922 14341 4924
rect 14397 4922 14421 4924
rect 14477 4922 14483 4924
rect 14237 4870 14239 4922
rect 14419 4870 14421 4922
rect 14175 4868 14181 4870
rect 14237 4868 14261 4870
rect 14317 4868 14341 4870
rect 14397 4868 14421 4870
rect 14477 4868 14483 4870
rect 14175 4859 14483 4868
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 12990 4176 13046 4185
rect 12990 4111 13046 4120
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12084 3126 12112 3470
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 11624 2854 11652 2994
rect 12176 2922 12204 3470
rect 12452 3194 12480 3674
rect 12912 3602 12940 3878
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12912 3058 12940 3538
rect 13004 3534 13032 4111
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13464 3534 13492 3878
rect 13648 3738 13676 4558
rect 13740 4486 13768 4762
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13740 4214 13768 4422
rect 14835 4380 15143 4389
rect 14835 4378 14841 4380
rect 14897 4378 14921 4380
rect 14977 4378 15001 4380
rect 15057 4378 15081 4380
rect 15137 4378 15143 4380
rect 14897 4326 14899 4378
rect 15079 4326 15081 4378
rect 14835 4324 14841 4326
rect 14897 4324 14921 4326
rect 14977 4324 15001 4326
rect 15057 4324 15081 4326
rect 15137 4324 15143 4326
rect 14835 4315 15143 4324
rect 15212 4282 15240 4626
rect 15396 4622 15424 4966
rect 15764 4826 15792 6718
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 16040 5914 16068 6190
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 16408 5234 16436 8230
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16684 7002 16712 7754
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16868 6798 16896 8910
rect 17420 8634 17448 8910
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17696 8090 17724 8366
rect 18616 8294 18644 9522
rect 19352 9450 19380 9930
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19465 9276 19773 9285
rect 19465 9274 19471 9276
rect 19527 9274 19551 9276
rect 19607 9274 19631 9276
rect 19687 9274 19711 9276
rect 19767 9274 19773 9276
rect 19527 9222 19529 9274
rect 19709 9222 19711 9274
rect 19465 9220 19471 9222
rect 19527 9220 19551 9222
rect 19607 9220 19631 9222
rect 19687 9220 19711 9222
rect 19767 9220 19773 9222
rect 19465 9211 19773 9220
rect 19996 9110 20024 12294
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20125 11996 20433 12005
rect 20125 11994 20131 11996
rect 20187 11994 20211 11996
rect 20267 11994 20291 11996
rect 20347 11994 20371 11996
rect 20427 11994 20433 11996
rect 20187 11942 20189 11994
rect 20369 11942 20371 11994
rect 20125 11940 20131 11942
rect 20187 11940 20211 11942
rect 20267 11940 20291 11942
rect 20347 11940 20371 11942
rect 20427 11940 20433 11942
rect 20125 11931 20433 11940
rect 20548 11898 20576 12038
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20640 11218 20668 12922
rect 20732 12442 20760 13262
rect 20720 12436 20772 12442
rect 20772 12406 20852 12434
rect 20720 12378 20772 12384
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20732 11898 20760 12174
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20125 10908 20433 10917
rect 20125 10906 20131 10908
rect 20187 10906 20211 10908
rect 20267 10906 20291 10908
rect 20347 10906 20371 10908
rect 20427 10906 20433 10908
rect 20187 10854 20189 10906
rect 20369 10854 20371 10906
rect 20125 10852 20131 10854
rect 20187 10852 20211 10854
rect 20267 10852 20291 10854
rect 20347 10852 20371 10854
rect 20427 10852 20433 10854
rect 20125 10843 20433 10852
rect 20548 10266 20576 11018
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20125 9820 20433 9829
rect 20125 9818 20131 9820
rect 20187 9818 20211 9820
rect 20267 9818 20291 9820
rect 20347 9818 20371 9820
rect 20427 9818 20433 9820
rect 20187 9766 20189 9818
rect 20369 9766 20371 9818
rect 20125 9764 20131 9766
rect 20187 9764 20211 9766
rect 20267 9764 20291 9766
rect 20347 9764 20371 9766
rect 20427 9764 20433 9766
rect 20125 9755 20433 9764
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20456 9178 20484 9522
rect 20548 9518 20576 9998
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 20548 9042 20576 9454
rect 20640 9450 20668 11018
rect 20732 10266 20760 11630
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20824 10146 20852 12406
rect 20996 12164 21048 12170
rect 20996 12106 21048 12112
rect 21008 11830 21036 12106
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21284 11354 21312 11698
rect 21376 11354 21404 13262
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21468 12442 21496 12582
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 22192 11688 22244 11694
rect 22190 11656 22192 11665
rect 22244 11656 22246 11665
rect 22190 11591 22246 11600
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 20732 10118 20852 10146
rect 20732 10062 20760 10118
rect 21008 10062 21036 10406
rect 21652 10266 21680 10406
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19904 8634 19932 8910
rect 20125 8732 20433 8741
rect 20125 8730 20131 8732
rect 20187 8730 20211 8732
rect 20267 8730 20291 8732
rect 20347 8730 20371 8732
rect 20427 8730 20433 8732
rect 20187 8678 20189 8730
rect 20369 8678 20371 8730
rect 20125 8676 20131 8678
rect 20187 8676 20211 8678
rect 20267 8676 20291 8678
rect 20347 8676 20371 8678
rect 20427 8676 20433 8678
rect 20125 8667 20433 8676
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16960 6798 16988 7142
rect 17512 6798 17540 7278
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 16868 6662 16896 6734
rect 17604 6730 17632 6938
rect 17696 6934 17724 8026
rect 18064 7954 18092 8230
rect 19465 8188 19773 8197
rect 19465 8186 19471 8188
rect 19527 8186 19551 8188
rect 19607 8186 19631 8188
rect 19687 8186 19711 8188
rect 19767 8186 19773 8188
rect 19527 8134 19529 8186
rect 19709 8134 19711 8186
rect 19465 8132 19471 8134
rect 19527 8132 19551 8134
rect 19607 8132 19631 8134
rect 19687 8132 19711 8134
rect 19767 8132 19773 8134
rect 19465 8123 19773 8132
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18064 7426 18092 7890
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 17972 7398 18092 7426
rect 17972 7002 18000 7398
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 7002 18092 7278
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 17684 6928 17736 6934
rect 17684 6870 17736 6876
rect 17696 6730 17724 6870
rect 17788 6866 17908 6882
rect 17788 6860 17920 6866
rect 17788 6854 17868 6860
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17684 6724 17736 6730
rect 17684 6666 17736 6672
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 16868 6118 16896 6598
rect 17420 6458 17448 6598
rect 17788 6458 17816 6854
rect 17868 6802 17920 6808
rect 18432 6798 18460 7686
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17880 6458 17908 6666
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16500 5914 16528 6054
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16868 5710 16896 6054
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 16040 4826 16068 5170
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16316 4826 16344 5102
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 15396 4282 15424 4558
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13740 3534 13768 4150
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14175 3836 14483 3845
rect 14175 3834 14181 3836
rect 14237 3834 14261 3836
rect 14317 3834 14341 3836
rect 14397 3834 14421 3836
rect 14477 3834 14483 3836
rect 14237 3782 14239 3834
rect 14419 3782 14421 3834
rect 14175 3780 14181 3782
rect 14237 3780 14261 3782
rect 14317 3780 14341 3782
rect 14397 3780 14421 3782
rect 14477 3780 14483 3782
rect 14175 3771 14483 3780
rect 12992 3528 13044 3534
rect 13176 3528 13228 3534
rect 12992 3470 13044 3476
rect 13096 3488 13176 3516
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 3595 2748 3903 2757
rect 3595 2746 3601 2748
rect 3657 2746 3681 2748
rect 3737 2746 3761 2748
rect 3817 2746 3841 2748
rect 3897 2746 3903 2748
rect 3657 2694 3659 2746
rect 3839 2694 3841 2746
rect 3595 2692 3601 2694
rect 3657 2692 3681 2694
rect 3737 2692 3761 2694
rect 3817 2692 3841 2694
rect 3897 2692 3903 2694
rect 3595 2683 3903 2692
rect 8588 2446 8616 2790
rect 8885 2748 9193 2757
rect 8885 2746 8891 2748
rect 8947 2746 8971 2748
rect 9027 2746 9051 2748
rect 9107 2746 9131 2748
rect 9187 2746 9193 2748
rect 8947 2694 8949 2746
rect 9129 2694 9131 2746
rect 8885 2692 8891 2694
rect 8947 2692 8971 2694
rect 9027 2692 9051 2694
rect 9107 2692 9131 2694
rect 9187 2692 9193 2694
rect 8885 2683 9193 2692
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 32 800 60 2382
rect 13096 2310 13124 3488
rect 13176 3470 13228 3476
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13188 2650 13216 2994
rect 13280 2854 13308 3334
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13464 2774 13492 3334
rect 14752 3194 14780 3878
rect 15672 3738 15700 4558
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16120 4208 16172 4214
rect 16120 4150 16172 4156
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 16132 3602 16160 4150
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 14835 3292 15143 3301
rect 14835 3290 14841 3292
rect 14897 3290 14921 3292
rect 14977 3290 15001 3292
rect 15057 3290 15081 3292
rect 15137 3290 15143 3292
rect 14897 3238 14899 3290
rect 15079 3238 15081 3290
rect 14835 3236 14841 3238
rect 14897 3236 14921 3238
rect 14977 3236 15001 3238
rect 15057 3236 15081 3238
rect 15137 3236 15143 3238
rect 14835 3227 15143 3236
rect 16224 3194 16252 4422
rect 16684 4282 16712 4558
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16500 3738 16528 4150
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16408 3194 16436 3538
rect 16592 3534 16620 3878
rect 16868 3738 16896 4490
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 17052 3534 17080 4150
rect 17144 3534 17172 5170
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17236 4826 17264 4966
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17880 4622 17908 6258
rect 18064 6118 18092 6598
rect 18800 6322 18828 6598
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 18064 5234 18092 5510
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16684 2990 16712 3402
rect 17144 3194 17172 3470
rect 17696 3346 17724 4218
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17788 3534 17816 3878
rect 17880 3738 17908 4218
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17880 3346 17908 3402
rect 17696 3318 17908 3346
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 13464 2746 13584 2774
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13556 2446 13584 2746
rect 14175 2748 14483 2757
rect 14175 2746 14181 2748
rect 14237 2746 14261 2748
rect 14317 2746 14341 2748
rect 14397 2746 14421 2748
rect 14477 2746 14483 2748
rect 14237 2694 14239 2746
rect 14419 2694 14421 2746
rect 14175 2692 14181 2694
rect 14237 2692 14261 2694
rect 14317 2692 14341 2694
rect 14397 2692 14421 2694
rect 14477 2692 14483 2694
rect 14175 2683 14483 2692
rect 17144 2514 17172 3130
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17512 2650 17540 2994
rect 17972 2650 18000 3606
rect 18064 3398 18092 4014
rect 18156 3942 18184 5646
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18432 4282 18460 4422
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18524 3738 18552 4558
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18708 4214 18736 4422
rect 18696 4208 18748 4214
rect 18696 4150 18748 4156
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18156 3194 18184 3470
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18524 2854 18552 3334
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18512 2848 18564 2854
rect 18512 2790 18564 2796
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 18524 2514 18552 2790
rect 18892 2650 18920 2994
rect 18984 2650 19012 7958
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 7410 19288 7686
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19352 7002 19380 7822
rect 20125 7644 20433 7653
rect 20125 7642 20131 7644
rect 20187 7642 20211 7644
rect 20267 7642 20291 7644
rect 20347 7642 20371 7644
rect 20427 7642 20433 7644
rect 20187 7590 20189 7642
rect 20369 7590 20371 7642
rect 20125 7588 20131 7590
rect 20187 7588 20211 7590
rect 20267 7588 20291 7590
rect 20347 7588 20371 7590
rect 20427 7588 20433 7590
rect 20125 7579 20433 7588
rect 20548 7478 20576 8978
rect 20732 8906 20760 9998
rect 20916 9654 20944 9998
rect 20904 9648 20956 9654
rect 20904 9590 20956 9596
rect 21008 9382 21036 9998
rect 21088 9988 21140 9994
rect 21088 9930 21140 9936
rect 21100 9722 21128 9930
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21284 9722 21312 9862
rect 21088 9716 21140 9722
rect 21272 9716 21324 9722
rect 21140 9676 21220 9704
rect 21088 9658 21140 9664
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21100 8974 21128 9318
rect 21192 9178 21220 9676
rect 21272 9658 21324 9664
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20732 7886 20760 8842
rect 21192 8498 21220 9114
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 20640 7546 20668 7822
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19465 7100 19773 7109
rect 19465 7098 19471 7100
rect 19527 7098 19551 7100
rect 19607 7098 19631 7100
rect 19687 7098 19711 7100
rect 19767 7098 19773 7100
rect 19527 7046 19529 7098
rect 19709 7046 19711 7098
rect 19465 7044 19471 7046
rect 19527 7044 19551 7046
rect 19607 7044 19631 7046
rect 19687 7044 19711 7046
rect 19767 7044 19773 7046
rect 19465 7035 19773 7044
rect 19904 7002 19932 7278
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 19904 6458 19932 6938
rect 19996 6730 20024 7414
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 20180 6662 20208 7346
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20456 6662 20484 7142
rect 20548 6866 20576 7414
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20125 6556 20433 6565
rect 20125 6554 20131 6556
rect 20187 6554 20211 6556
rect 20267 6554 20291 6556
rect 20347 6554 20371 6556
rect 20427 6554 20433 6556
rect 20187 6502 20189 6554
rect 20369 6502 20371 6554
rect 20125 6500 20131 6502
rect 20187 6500 20211 6502
rect 20267 6500 20291 6502
rect 20347 6500 20371 6502
rect 20427 6500 20433 6502
rect 20125 6491 20433 6500
rect 19892 6452 19944 6458
rect 19892 6394 19944 6400
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19352 5370 19380 6054
rect 19465 6012 19773 6021
rect 19465 6010 19471 6012
rect 19527 6010 19551 6012
rect 19607 6010 19631 6012
rect 19687 6010 19711 6012
rect 19767 6010 19773 6012
rect 19527 5958 19529 6010
rect 19709 5958 19711 6010
rect 19465 5956 19471 5958
rect 19527 5956 19551 5958
rect 19607 5956 19631 5958
rect 19687 5956 19711 5958
rect 19767 5956 19773 5958
rect 19465 5947 19773 5956
rect 19904 5778 19932 6394
rect 20548 6390 20576 6802
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 19892 5568 19944 5574
rect 19892 5510 19944 5516
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19904 5234 19932 5510
rect 19996 5370 20024 6326
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20272 5914 20300 6258
rect 20640 6118 20668 7346
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20125 5468 20433 5477
rect 20125 5466 20131 5468
rect 20187 5466 20211 5468
rect 20267 5466 20291 5468
rect 20347 5466 20371 5468
rect 20427 5466 20433 5468
rect 20187 5414 20189 5466
rect 20369 5414 20371 5466
rect 20125 5412 20131 5414
rect 20187 5412 20211 5414
rect 20267 5412 20291 5414
rect 20347 5412 20371 5414
rect 20427 5412 20433 5414
rect 20125 5403 20433 5412
rect 20548 5370 20576 5646
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19465 4924 19773 4933
rect 19465 4922 19471 4924
rect 19527 4922 19551 4924
rect 19607 4922 19631 4924
rect 19687 4922 19711 4924
rect 19767 4922 19773 4924
rect 19527 4870 19529 4922
rect 19709 4870 19711 4922
rect 19465 4868 19471 4870
rect 19527 4868 19551 4870
rect 19607 4868 19631 4870
rect 19687 4868 19711 4870
rect 19767 4868 19773 4870
rect 19465 4859 19773 4868
rect 19996 4282 20024 5306
rect 20640 5234 20668 5510
rect 20732 5370 20760 7822
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 20824 6798 20852 7686
rect 21560 7410 21588 7686
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21192 5778 21220 6054
rect 21180 5772 21232 5778
rect 21180 5714 21232 5720
rect 21836 5370 21864 7822
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20125 4380 20433 4389
rect 20125 4378 20131 4380
rect 20187 4378 20211 4380
rect 20267 4378 20291 4380
rect 20347 4378 20371 4380
rect 20427 4378 20433 4380
rect 20187 4326 20189 4378
rect 20369 4326 20371 4378
rect 20125 4324 20131 4326
rect 20187 4324 20211 4326
rect 20267 4324 20291 4326
rect 20347 4324 20371 4326
rect 20427 4324 20433 4326
rect 20125 4315 20433 4324
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 19352 3194 19380 4082
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19465 3836 19773 3845
rect 19465 3834 19471 3836
rect 19527 3834 19551 3836
rect 19607 3834 19631 3836
rect 19687 3834 19711 3836
rect 19767 3834 19773 3836
rect 19527 3782 19529 3834
rect 19709 3782 19711 3834
rect 19465 3780 19471 3782
rect 19527 3780 19551 3782
rect 19607 3780 19631 3782
rect 19687 3780 19711 3782
rect 19767 3780 19773 3782
rect 19465 3771 19773 3780
rect 19812 3534 19840 3878
rect 20180 3738 20208 4082
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 19996 3194 20024 3470
rect 20125 3292 20433 3301
rect 20125 3290 20131 3292
rect 20187 3290 20211 3292
rect 20267 3290 20291 3292
rect 20347 3290 20371 3292
rect 20427 3290 20433 3292
rect 20187 3238 20189 3290
rect 20369 3238 20371 3290
rect 20125 3236 20131 3238
rect 20187 3236 20211 3238
rect 20267 3236 20291 3238
rect 20347 3236 20371 3238
rect 20427 3236 20433 3238
rect 20125 3227 20433 3236
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 19465 2748 19773 2757
rect 19465 2746 19471 2748
rect 19527 2746 19551 2748
rect 19607 2746 19631 2748
rect 19687 2746 19711 2748
rect 19767 2746 19773 2748
rect 19527 2694 19529 2746
rect 19709 2694 19711 2746
rect 19465 2692 19471 2694
rect 19527 2692 19551 2694
rect 19607 2692 19631 2694
rect 19687 2692 19711 2694
rect 19767 2692 19773 2694
rect 19465 2683 19773 2692
rect 21468 2650 21496 2994
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 18512 2508 18564 2514
rect 18512 2450 18564 2456
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 17868 2372 17920 2378
rect 17868 2314 17920 2320
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 4255 2204 4563 2213
rect 4255 2202 4261 2204
rect 4317 2202 4341 2204
rect 4397 2202 4421 2204
rect 4477 2202 4501 2204
rect 4557 2202 4563 2204
rect 4317 2150 4319 2202
rect 4499 2150 4501 2202
rect 4255 2148 4261 2150
rect 4317 2148 4341 2150
rect 4397 2148 4421 2150
rect 4477 2148 4501 2150
rect 4557 2148 4563 2150
rect 4255 2139 4563 2148
rect 8404 800 8432 2246
rect 9545 2204 9853 2213
rect 9545 2202 9551 2204
rect 9607 2202 9631 2204
rect 9687 2202 9711 2204
rect 9767 2202 9791 2204
rect 9847 2202 9853 2204
rect 9607 2150 9609 2202
rect 9789 2150 9791 2202
rect 9545 2148 9551 2150
rect 9607 2148 9631 2150
rect 9687 2148 9711 2150
rect 9767 2148 9791 2150
rect 9847 2148 9853 2150
rect 9545 2139 9853 2148
rect 14835 2204 15143 2213
rect 14835 2202 14841 2204
rect 14897 2202 14921 2204
rect 14977 2202 15001 2204
rect 15057 2202 15081 2204
rect 15137 2202 15143 2204
rect 14897 2150 14899 2202
rect 15079 2150 15081 2202
rect 14835 2148 14841 2150
rect 14897 2148 14921 2150
rect 14977 2148 15001 2150
rect 15057 2148 15081 2150
rect 15137 2148 15143 2150
rect 14835 2139 15143 2148
rect 17420 870 17540 898
rect 17420 800 17448 870
rect 18 0 74 800
rect 8390 0 8446 800
rect 17406 0 17462 800
rect 17512 762 17540 870
rect 17880 762 17908 2314
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 20125 2204 20433 2213
rect 20125 2202 20131 2204
rect 20187 2202 20211 2204
rect 20267 2202 20291 2204
rect 20347 2202 20371 2204
rect 20427 2202 20433 2204
rect 20187 2150 20189 2202
rect 20369 2150 20371 2202
rect 20125 2148 20131 2150
rect 20187 2148 20211 2150
rect 20267 2148 20291 2150
rect 20347 2148 20371 2150
rect 20427 2148 20433 2150
rect 20125 2139 20433 2148
rect 22204 2145 22232 2246
rect 22190 2136 22246 2145
rect 22190 2071 22246 2080
rect 17512 734 17908 762
<< via2 >>
rect 4261 22874 4317 22876
rect 4341 22874 4397 22876
rect 4421 22874 4477 22876
rect 4501 22874 4557 22876
rect 4261 22822 4307 22874
rect 4307 22822 4317 22874
rect 4341 22822 4371 22874
rect 4371 22822 4383 22874
rect 4383 22822 4397 22874
rect 4421 22822 4435 22874
rect 4435 22822 4447 22874
rect 4447 22822 4477 22874
rect 4501 22822 4511 22874
rect 4511 22822 4557 22874
rect 4261 22820 4317 22822
rect 4341 22820 4397 22822
rect 4421 22820 4477 22822
rect 4501 22820 4557 22822
rect 9551 22874 9607 22876
rect 9631 22874 9687 22876
rect 9711 22874 9767 22876
rect 9791 22874 9847 22876
rect 9551 22822 9597 22874
rect 9597 22822 9607 22874
rect 9631 22822 9661 22874
rect 9661 22822 9673 22874
rect 9673 22822 9687 22874
rect 9711 22822 9725 22874
rect 9725 22822 9737 22874
rect 9737 22822 9767 22874
rect 9791 22822 9801 22874
rect 9801 22822 9847 22874
rect 9551 22820 9607 22822
rect 9631 22820 9687 22822
rect 9711 22820 9767 22822
rect 9791 22820 9847 22822
rect 14841 22874 14897 22876
rect 14921 22874 14977 22876
rect 15001 22874 15057 22876
rect 15081 22874 15137 22876
rect 14841 22822 14887 22874
rect 14887 22822 14897 22874
rect 14921 22822 14951 22874
rect 14951 22822 14963 22874
rect 14963 22822 14977 22874
rect 15001 22822 15015 22874
rect 15015 22822 15027 22874
rect 15027 22822 15057 22874
rect 15081 22822 15091 22874
rect 15091 22822 15137 22874
rect 14841 22820 14897 22822
rect 14921 22820 14977 22822
rect 15001 22820 15057 22822
rect 15081 22820 15137 22822
rect 20131 22874 20187 22876
rect 20211 22874 20267 22876
rect 20291 22874 20347 22876
rect 20371 22874 20427 22876
rect 20131 22822 20177 22874
rect 20177 22822 20187 22874
rect 20211 22822 20241 22874
rect 20241 22822 20253 22874
rect 20253 22822 20267 22874
rect 20291 22822 20305 22874
rect 20305 22822 20317 22874
rect 20317 22822 20347 22874
rect 20371 22822 20381 22874
rect 20381 22822 20427 22874
rect 20131 22820 20187 22822
rect 20211 22820 20267 22822
rect 20291 22820 20347 22822
rect 20371 22820 20427 22822
rect 3601 22330 3657 22332
rect 3681 22330 3737 22332
rect 3761 22330 3817 22332
rect 3841 22330 3897 22332
rect 3601 22278 3647 22330
rect 3647 22278 3657 22330
rect 3681 22278 3711 22330
rect 3711 22278 3723 22330
rect 3723 22278 3737 22330
rect 3761 22278 3775 22330
rect 3775 22278 3787 22330
rect 3787 22278 3817 22330
rect 3841 22278 3851 22330
rect 3851 22278 3897 22330
rect 3601 22276 3657 22278
rect 3681 22276 3737 22278
rect 3761 22276 3817 22278
rect 3841 22276 3897 22278
rect 8891 22330 8947 22332
rect 8971 22330 9027 22332
rect 9051 22330 9107 22332
rect 9131 22330 9187 22332
rect 8891 22278 8937 22330
rect 8937 22278 8947 22330
rect 8971 22278 9001 22330
rect 9001 22278 9013 22330
rect 9013 22278 9027 22330
rect 9051 22278 9065 22330
rect 9065 22278 9077 22330
rect 9077 22278 9107 22330
rect 9131 22278 9141 22330
rect 9141 22278 9187 22330
rect 8891 22276 8947 22278
rect 8971 22276 9027 22278
rect 9051 22276 9107 22278
rect 9131 22276 9187 22278
rect 4261 21786 4317 21788
rect 4341 21786 4397 21788
rect 4421 21786 4477 21788
rect 4501 21786 4557 21788
rect 4261 21734 4307 21786
rect 4307 21734 4317 21786
rect 4341 21734 4371 21786
rect 4371 21734 4383 21786
rect 4383 21734 4397 21786
rect 4421 21734 4435 21786
rect 4435 21734 4447 21786
rect 4447 21734 4477 21786
rect 4501 21734 4511 21786
rect 4511 21734 4557 21786
rect 4261 21732 4317 21734
rect 4341 21732 4397 21734
rect 4421 21732 4477 21734
rect 4501 21732 4557 21734
rect 3601 21242 3657 21244
rect 3681 21242 3737 21244
rect 3761 21242 3817 21244
rect 3841 21242 3897 21244
rect 3601 21190 3647 21242
rect 3647 21190 3657 21242
rect 3681 21190 3711 21242
rect 3711 21190 3723 21242
rect 3723 21190 3737 21242
rect 3761 21190 3775 21242
rect 3775 21190 3787 21242
rect 3787 21190 3817 21242
rect 3841 21190 3851 21242
rect 3851 21190 3897 21242
rect 3601 21188 3657 21190
rect 3681 21188 3737 21190
rect 3761 21188 3817 21190
rect 3841 21188 3897 21190
rect 3601 20154 3657 20156
rect 3681 20154 3737 20156
rect 3761 20154 3817 20156
rect 3841 20154 3897 20156
rect 3601 20102 3647 20154
rect 3647 20102 3657 20154
rect 3681 20102 3711 20154
rect 3711 20102 3723 20154
rect 3723 20102 3737 20154
rect 3761 20102 3775 20154
rect 3775 20102 3787 20154
rect 3787 20102 3817 20154
rect 3841 20102 3851 20154
rect 3851 20102 3897 20154
rect 3601 20100 3657 20102
rect 3681 20100 3737 20102
rect 3761 20100 3817 20102
rect 3841 20100 3897 20102
rect 3601 19066 3657 19068
rect 3681 19066 3737 19068
rect 3761 19066 3817 19068
rect 3841 19066 3897 19068
rect 3601 19014 3647 19066
rect 3647 19014 3657 19066
rect 3681 19014 3711 19066
rect 3711 19014 3723 19066
rect 3723 19014 3737 19066
rect 3761 19014 3775 19066
rect 3775 19014 3787 19066
rect 3787 19014 3817 19066
rect 3841 19014 3851 19066
rect 3851 19014 3897 19066
rect 3601 19012 3657 19014
rect 3681 19012 3737 19014
rect 3761 19012 3817 19014
rect 3841 19012 3897 19014
rect 4261 20698 4317 20700
rect 4341 20698 4397 20700
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4261 20646 4307 20698
rect 4307 20646 4317 20698
rect 4341 20646 4371 20698
rect 4371 20646 4383 20698
rect 4383 20646 4397 20698
rect 4421 20646 4435 20698
rect 4435 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4261 20644 4317 20646
rect 4341 20644 4397 20646
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4261 19610 4317 19612
rect 4341 19610 4397 19612
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4261 19558 4307 19610
rect 4307 19558 4317 19610
rect 4341 19558 4371 19610
rect 4371 19558 4383 19610
rect 4383 19558 4397 19610
rect 4421 19558 4435 19610
rect 4435 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4261 19556 4317 19558
rect 4341 19556 4397 19558
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4261 18522 4317 18524
rect 4341 18522 4397 18524
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4261 18470 4307 18522
rect 4307 18470 4317 18522
rect 4341 18470 4371 18522
rect 4371 18470 4383 18522
rect 4383 18470 4397 18522
rect 4421 18470 4435 18522
rect 4435 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4261 18468 4317 18470
rect 4341 18468 4397 18470
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 3601 17978 3657 17980
rect 3681 17978 3737 17980
rect 3761 17978 3817 17980
rect 3841 17978 3897 17980
rect 3601 17926 3647 17978
rect 3647 17926 3657 17978
rect 3681 17926 3711 17978
rect 3711 17926 3723 17978
rect 3723 17926 3737 17978
rect 3761 17926 3775 17978
rect 3775 17926 3787 17978
rect 3787 17926 3817 17978
rect 3841 17926 3851 17978
rect 3851 17926 3897 17978
rect 3601 17924 3657 17926
rect 3681 17924 3737 17926
rect 3761 17924 3817 17926
rect 3841 17924 3897 17926
rect 4261 17434 4317 17436
rect 4341 17434 4397 17436
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4261 17382 4307 17434
rect 4307 17382 4317 17434
rect 4341 17382 4371 17434
rect 4371 17382 4383 17434
rect 4383 17382 4397 17434
rect 4421 17382 4435 17434
rect 4435 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4261 17380 4317 17382
rect 4341 17380 4397 17382
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 6734 21392 6790 21448
rect 7654 21392 7710 21448
rect 9551 21786 9607 21788
rect 9631 21786 9687 21788
rect 9711 21786 9767 21788
rect 9791 21786 9847 21788
rect 9551 21734 9597 21786
rect 9597 21734 9607 21786
rect 9631 21734 9661 21786
rect 9661 21734 9673 21786
rect 9673 21734 9687 21786
rect 9711 21734 9725 21786
rect 9725 21734 9737 21786
rect 9737 21734 9767 21786
rect 9791 21734 9801 21786
rect 9801 21734 9847 21786
rect 9551 21732 9607 21734
rect 9631 21732 9687 21734
rect 9711 21732 9767 21734
rect 9791 21732 9847 21734
rect 8891 21242 8947 21244
rect 8971 21242 9027 21244
rect 9051 21242 9107 21244
rect 9131 21242 9187 21244
rect 8891 21190 8937 21242
rect 8937 21190 8947 21242
rect 8971 21190 9001 21242
rect 9001 21190 9013 21242
rect 9013 21190 9027 21242
rect 9051 21190 9065 21242
rect 9065 21190 9077 21242
rect 9077 21190 9107 21242
rect 9131 21190 9141 21242
rect 9141 21190 9187 21242
rect 8891 21188 8947 21190
rect 8971 21188 9027 21190
rect 9051 21188 9107 21190
rect 9131 21188 9187 21190
rect 3601 16890 3657 16892
rect 3681 16890 3737 16892
rect 3761 16890 3817 16892
rect 3841 16890 3897 16892
rect 3601 16838 3647 16890
rect 3647 16838 3657 16890
rect 3681 16838 3711 16890
rect 3711 16838 3723 16890
rect 3723 16838 3737 16890
rect 3761 16838 3775 16890
rect 3775 16838 3787 16890
rect 3787 16838 3817 16890
rect 3841 16838 3851 16890
rect 3851 16838 3897 16890
rect 3601 16836 3657 16838
rect 3681 16836 3737 16838
rect 3761 16836 3817 16838
rect 3841 16836 3897 16838
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 4261 16346 4317 16348
rect 4341 16346 4397 16348
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4261 16294 4307 16346
rect 4307 16294 4317 16346
rect 4341 16294 4371 16346
rect 4371 16294 4383 16346
rect 4383 16294 4397 16346
rect 4421 16294 4435 16346
rect 4435 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4261 16292 4317 16294
rect 4341 16292 4397 16294
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 3601 15802 3657 15804
rect 3681 15802 3737 15804
rect 3761 15802 3817 15804
rect 3841 15802 3897 15804
rect 3601 15750 3647 15802
rect 3647 15750 3657 15802
rect 3681 15750 3711 15802
rect 3711 15750 3723 15802
rect 3723 15750 3737 15802
rect 3761 15750 3775 15802
rect 3775 15750 3787 15802
rect 3787 15750 3817 15802
rect 3841 15750 3851 15802
rect 3851 15750 3897 15802
rect 3601 15748 3657 15750
rect 3681 15748 3737 15750
rect 3761 15748 3817 15750
rect 3841 15748 3897 15750
rect 5078 18400 5134 18456
rect 4261 15258 4317 15260
rect 4341 15258 4397 15260
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4261 15206 4307 15258
rect 4307 15206 4317 15258
rect 4341 15206 4371 15258
rect 4371 15206 4383 15258
rect 4383 15206 4397 15258
rect 4421 15206 4435 15258
rect 4435 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4261 15204 4317 15206
rect 4341 15204 4397 15206
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 3601 14714 3657 14716
rect 3681 14714 3737 14716
rect 3761 14714 3817 14716
rect 3841 14714 3897 14716
rect 3601 14662 3647 14714
rect 3647 14662 3657 14714
rect 3681 14662 3711 14714
rect 3711 14662 3723 14714
rect 3723 14662 3737 14714
rect 3761 14662 3775 14714
rect 3775 14662 3787 14714
rect 3787 14662 3817 14714
rect 3841 14662 3851 14714
rect 3851 14662 3897 14714
rect 3601 14660 3657 14662
rect 3681 14660 3737 14662
rect 3761 14660 3817 14662
rect 3841 14660 3897 14662
rect 4261 14170 4317 14172
rect 4341 14170 4397 14172
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4261 14118 4307 14170
rect 4307 14118 4317 14170
rect 4341 14118 4371 14170
rect 4371 14118 4383 14170
rect 4383 14118 4397 14170
rect 4421 14118 4435 14170
rect 4435 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4261 14116 4317 14118
rect 4341 14116 4397 14118
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 3601 13626 3657 13628
rect 3681 13626 3737 13628
rect 3761 13626 3817 13628
rect 3841 13626 3897 13628
rect 3601 13574 3647 13626
rect 3647 13574 3657 13626
rect 3681 13574 3711 13626
rect 3711 13574 3723 13626
rect 3723 13574 3737 13626
rect 3761 13574 3775 13626
rect 3775 13574 3787 13626
rect 3787 13574 3817 13626
rect 3841 13574 3851 13626
rect 3851 13574 3897 13626
rect 3601 13572 3657 13574
rect 3681 13572 3737 13574
rect 3761 13572 3817 13574
rect 3841 13572 3897 13574
rect 3601 12538 3657 12540
rect 3681 12538 3737 12540
rect 3761 12538 3817 12540
rect 3841 12538 3897 12540
rect 3601 12486 3647 12538
rect 3647 12486 3657 12538
rect 3681 12486 3711 12538
rect 3711 12486 3723 12538
rect 3723 12486 3737 12538
rect 3761 12486 3775 12538
rect 3775 12486 3787 12538
rect 3787 12486 3817 12538
rect 3841 12486 3851 12538
rect 3851 12486 3897 12538
rect 3601 12484 3657 12486
rect 3681 12484 3737 12486
rect 3761 12484 3817 12486
rect 3841 12484 3897 12486
rect 4261 13082 4317 13084
rect 4341 13082 4397 13084
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4261 13030 4307 13082
rect 4307 13030 4317 13082
rect 4341 13030 4371 13082
rect 4371 13030 4383 13082
rect 4383 13030 4397 13082
rect 4421 13030 4435 13082
rect 4435 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4261 13028 4317 13030
rect 4341 13028 4397 13030
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4261 11994 4317 11996
rect 4341 11994 4397 11996
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4261 11942 4307 11994
rect 4307 11942 4317 11994
rect 4341 11942 4371 11994
rect 4371 11942 4383 11994
rect 4383 11942 4397 11994
rect 4421 11942 4435 11994
rect 4435 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4261 11940 4317 11942
rect 4341 11940 4397 11942
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 3601 11450 3657 11452
rect 3681 11450 3737 11452
rect 3761 11450 3817 11452
rect 3841 11450 3897 11452
rect 3601 11398 3647 11450
rect 3647 11398 3657 11450
rect 3681 11398 3711 11450
rect 3711 11398 3723 11450
rect 3723 11398 3737 11450
rect 3761 11398 3775 11450
rect 3775 11398 3787 11450
rect 3787 11398 3817 11450
rect 3841 11398 3851 11450
rect 3851 11398 3897 11450
rect 3601 11396 3657 11398
rect 3681 11396 3737 11398
rect 3761 11396 3817 11398
rect 3841 11396 3897 11398
rect 4261 10906 4317 10908
rect 4341 10906 4397 10908
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4261 10854 4307 10906
rect 4307 10854 4317 10906
rect 4341 10854 4371 10906
rect 4371 10854 4383 10906
rect 4383 10854 4397 10906
rect 4421 10854 4435 10906
rect 4435 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4261 10852 4317 10854
rect 4341 10852 4397 10854
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 3601 10362 3657 10364
rect 3681 10362 3737 10364
rect 3761 10362 3817 10364
rect 3841 10362 3897 10364
rect 3601 10310 3647 10362
rect 3647 10310 3657 10362
rect 3681 10310 3711 10362
rect 3711 10310 3723 10362
rect 3723 10310 3737 10362
rect 3761 10310 3775 10362
rect 3775 10310 3787 10362
rect 3787 10310 3817 10362
rect 3841 10310 3851 10362
rect 3851 10310 3897 10362
rect 3601 10308 3657 10310
rect 3681 10308 3737 10310
rect 3761 10308 3817 10310
rect 3841 10308 3897 10310
rect 4261 9818 4317 9820
rect 4341 9818 4397 9820
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4261 9766 4307 9818
rect 4307 9766 4317 9818
rect 4341 9766 4371 9818
rect 4371 9766 4383 9818
rect 4383 9766 4397 9818
rect 4421 9766 4435 9818
rect 4435 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4261 9764 4317 9766
rect 4341 9764 4397 9766
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 3601 9274 3657 9276
rect 3681 9274 3737 9276
rect 3761 9274 3817 9276
rect 3841 9274 3897 9276
rect 3601 9222 3647 9274
rect 3647 9222 3657 9274
rect 3681 9222 3711 9274
rect 3711 9222 3723 9274
rect 3723 9222 3737 9274
rect 3761 9222 3775 9274
rect 3775 9222 3787 9274
rect 3787 9222 3817 9274
rect 3841 9222 3851 9274
rect 3851 9222 3897 9274
rect 3601 9220 3657 9222
rect 3681 9220 3737 9222
rect 3761 9220 3817 9222
rect 3841 9220 3897 9222
rect 3601 8186 3657 8188
rect 3681 8186 3737 8188
rect 3761 8186 3817 8188
rect 3841 8186 3897 8188
rect 3601 8134 3647 8186
rect 3647 8134 3657 8186
rect 3681 8134 3711 8186
rect 3711 8134 3723 8186
rect 3723 8134 3737 8186
rect 3761 8134 3775 8186
rect 3775 8134 3787 8186
rect 3787 8134 3817 8186
rect 3841 8134 3851 8186
rect 3851 8134 3897 8186
rect 3601 8132 3657 8134
rect 3681 8132 3737 8134
rect 3761 8132 3817 8134
rect 3841 8132 3897 8134
rect 3601 7098 3657 7100
rect 3681 7098 3737 7100
rect 3761 7098 3817 7100
rect 3841 7098 3897 7100
rect 3601 7046 3647 7098
rect 3647 7046 3657 7098
rect 3681 7046 3711 7098
rect 3711 7046 3723 7098
rect 3723 7046 3737 7098
rect 3761 7046 3775 7098
rect 3775 7046 3787 7098
rect 3787 7046 3817 7098
rect 3841 7046 3851 7098
rect 3851 7046 3897 7098
rect 3601 7044 3657 7046
rect 3681 7044 3737 7046
rect 3761 7044 3817 7046
rect 3841 7044 3897 7046
rect 3601 6010 3657 6012
rect 3681 6010 3737 6012
rect 3761 6010 3817 6012
rect 3841 6010 3897 6012
rect 3601 5958 3647 6010
rect 3647 5958 3657 6010
rect 3681 5958 3711 6010
rect 3711 5958 3723 6010
rect 3723 5958 3737 6010
rect 3761 5958 3775 6010
rect 3775 5958 3787 6010
rect 3787 5958 3817 6010
rect 3841 5958 3851 6010
rect 3851 5958 3897 6010
rect 3601 5956 3657 5958
rect 3681 5956 3737 5958
rect 3761 5956 3817 5958
rect 3841 5956 3897 5958
rect 4261 8730 4317 8732
rect 4341 8730 4397 8732
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4261 8678 4307 8730
rect 4307 8678 4317 8730
rect 4341 8678 4371 8730
rect 4371 8678 4383 8730
rect 4383 8678 4397 8730
rect 4421 8678 4435 8730
rect 4435 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4261 8676 4317 8678
rect 4341 8676 4397 8678
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4261 7642 4317 7644
rect 4341 7642 4397 7644
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4261 7590 4307 7642
rect 4307 7590 4317 7642
rect 4341 7590 4371 7642
rect 4371 7590 4383 7642
rect 4383 7590 4397 7642
rect 4421 7590 4435 7642
rect 4435 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4261 7588 4317 7590
rect 4341 7588 4397 7590
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 8891 20154 8947 20156
rect 8971 20154 9027 20156
rect 9051 20154 9107 20156
rect 9131 20154 9187 20156
rect 8891 20102 8937 20154
rect 8937 20102 8947 20154
rect 8971 20102 9001 20154
rect 9001 20102 9013 20154
rect 9013 20102 9027 20154
rect 9051 20102 9065 20154
rect 9065 20102 9077 20154
rect 9077 20102 9107 20154
rect 9131 20102 9141 20154
rect 9141 20102 9187 20154
rect 8891 20100 8947 20102
rect 8971 20100 9027 20102
rect 9051 20100 9107 20102
rect 9131 20100 9187 20102
rect 8891 19066 8947 19068
rect 8971 19066 9027 19068
rect 9051 19066 9107 19068
rect 9131 19066 9187 19068
rect 8891 19014 8937 19066
rect 8937 19014 8947 19066
rect 8971 19014 9001 19066
rect 9001 19014 9013 19066
rect 9013 19014 9027 19066
rect 9051 19014 9065 19066
rect 9065 19014 9077 19066
rect 9077 19014 9107 19066
rect 9131 19014 9141 19066
rect 9141 19014 9187 19066
rect 8891 19012 8947 19014
rect 8971 19012 9027 19014
rect 9051 19012 9107 19014
rect 9131 19012 9187 19014
rect 8891 17978 8947 17980
rect 8971 17978 9027 17980
rect 9051 17978 9107 17980
rect 9131 17978 9187 17980
rect 8891 17926 8937 17978
rect 8937 17926 8947 17978
rect 8971 17926 9001 17978
rect 9001 17926 9013 17978
rect 9013 17926 9027 17978
rect 9051 17926 9065 17978
rect 9065 17926 9077 17978
rect 9077 17926 9107 17978
rect 9131 17926 9141 17978
rect 9141 17926 9187 17978
rect 8891 17924 8947 17926
rect 8971 17924 9027 17926
rect 9051 17924 9107 17926
rect 9131 17924 9187 17926
rect 9551 20698 9607 20700
rect 9631 20698 9687 20700
rect 9711 20698 9767 20700
rect 9791 20698 9847 20700
rect 9551 20646 9597 20698
rect 9597 20646 9607 20698
rect 9631 20646 9661 20698
rect 9661 20646 9673 20698
rect 9673 20646 9687 20698
rect 9711 20646 9725 20698
rect 9725 20646 9737 20698
rect 9737 20646 9767 20698
rect 9791 20646 9801 20698
rect 9801 20646 9847 20698
rect 9551 20644 9607 20646
rect 9631 20644 9687 20646
rect 9711 20644 9767 20646
rect 9791 20644 9847 20646
rect 9551 19610 9607 19612
rect 9631 19610 9687 19612
rect 9711 19610 9767 19612
rect 9791 19610 9847 19612
rect 9551 19558 9597 19610
rect 9597 19558 9607 19610
rect 9631 19558 9661 19610
rect 9661 19558 9673 19610
rect 9673 19558 9687 19610
rect 9711 19558 9725 19610
rect 9725 19558 9737 19610
rect 9737 19558 9767 19610
rect 9791 19558 9801 19610
rect 9801 19558 9847 19610
rect 9551 19556 9607 19558
rect 9631 19556 9687 19558
rect 9711 19556 9767 19558
rect 9791 19556 9847 19558
rect 11334 19352 11390 19408
rect 12162 19352 12218 19408
rect 9551 18522 9607 18524
rect 9631 18522 9687 18524
rect 9711 18522 9767 18524
rect 9791 18522 9847 18524
rect 9551 18470 9597 18522
rect 9597 18470 9607 18522
rect 9631 18470 9661 18522
rect 9661 18470 9673 18522
rect 9673 18470 9687 18522
rect 9711 18470 9725 18522
rect 9725 18470 9737 18522
rect 9737 18470 9767 18522
rect 9791 18470 9801 18522
rect 9801 18470 9847 18522
rect 9551 18468 9607 18470
rect 9631 18468 9687 18470
rect 9711 18468 9767 18470
rect 9791 18468 9847 18470
rect 9218 17176 9274 17232
rect 9551 17434 9607 17436
rect 9631 17434 9687 17436
rect 9711 17434 9767 17436
rect 9791 17434 9847 17436
rect 9551 17382 9597 17434
rect 9597 17382 9607 17434
rect 9631 17382 9661 17434
rect 9661 17382 9673 17434
rect 9673 17382 9687 17434
rect 9711 17382 9725 17434
rect 9725 17382 9737 17434
rect 9737 17382 9767 17434
rect 9791 17382 9801 17434
rect 9801 17382 9847 17434
rect 9551 17380 9607 17382
rect 9631 17380 9687 17382
rect 9711 17380 9767 17382
rect 9791 17380 9847 17382
rect 9494 17212 9496 17232
rect 9496 17212 9548 17232
rect 9548 17212 9550 17232
rect 9494 17176 9550 17212
rect 8891 16890 8947 16892
rect 8971 16890 9027 16892
rect 9051 16890 9107 16892
rect 9131 16890 9187 16892
rect 8891 16838 8937 16890
rect 8937 16838 8947 16890
rect 8971 16838 9001 16890
rect 9001 16838 9013 16890
rect 9013 16838 9027 16890
rect 9051 16838 9065 16890
rect 9065 16838 9077 16890
rect 9077 16838 9107 16890
rect 9131 16838 9141 16890
rect 9141 16838 9187 16890
rect 8891 16836 8947 16838
rect 8971 16836 9027 16838
rect 9051 16836 9107 16838
rect 9131 16836 9187 16838
rect 9551 16346 9607 16348
rect 9631 16346 9687 16348
rect 9711 16346 9767 16348
rect 9791 16346 9847 16348
rect 9551 16294 9597 16346
rect 9597 16294 9607 16346
rect 9631 16294 9661 16346
rect 9661 16294 9673 16346
rect 9673 16294 9687 16346
rect 9711 16294 9725 16346
rect 9725 16294 9737 16346
rect 9737 16294 9767 16346
rect 9791 16294 9801 16346
rect 9801 16294 9847 16346
rect 9551 16292 9607 16294
rect 9631 16292 9687 16294
rect 9711 16292 9767 16294
rect 9791 16292 9847 16294
rect 8891 15802 8947 15804
rect 8971 15802 9027 15804
rect 9051 15802 9107 15804
rect 9131 15802 9187 15804
rect 8891 15750 8937 15802
rect 8937 15750 8947 15802
rect 8971 15750 9001 15802
rect 9001 15750 9013 15802
rect 9013 15750 9027 15802
rect 9051 15750 9065 15802
rect 9065 15750 9077 15802
rect 9077 15750 9107 15802
rect 9131 15750 9141 15802
rect 9141 15750 9187 15802
rect 8891 15748 8947 15750
rect 8971 15748 9027 15750
rect 9051 15748 9107 15750
rect 9131 15748 9187 15750
rect 9551 15258 9607 15260
rect 9631 15258 9687 15260
rect 9711 15258 9767 15260
rect 9791 15258 9847 15260
rect 9551 15206 9597 15258
rect 9597 15206 9607 15258
rect 9631 15206 9661 15258
rect 9661 15206 9673 15258
rect 9673 15206 9687 15258
rect 9711 15206 9725 15258
rect 9725 15206 9737 15258
rect 9737 15206 9767 15258
rect 9791 15206 9801 15258
rect 9801 15206 9847 15258
rect 9551 15204 9607 15206
rect 9631 15204 9687 15206
rect 9711 15204 9767 15206
rect 9791 15204 9847 15206
rect 8891 14714 8947 14716
rect 8971 14714 9027 14716
rect 9051 14714 9107 14716
rect 9131 14714 9187 14716
rect 8891 14662 8937 14714
rect 8937 14662 8947 14714
rect 8971 14662 9001 14714
rect 9001 14662 9013 14714
rect 9013 14662 9027 14714
rect 9051 14662 9065 14714
rect 9065 14662 9077 14714
rect 9077 14662 9107 14714
rect 9131 14662 9141 14714
rect 9141 14662 9187 14714
rect 8891 14660 8947 14662
rect 8971 14660 9027 14662
rect 9051 14660 9107 14662
rect 9131 14660 9187 14662
rect 4261 6554 4317 6556
rect 4341 6554 4397 6556
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4261 6502 4307 6554
rect 4307 6502 4317 6554
rect 4341 6502 4371 6554
rect 4371 6502 4383 6554
rect 4383 6502 4397 6554
rect 4421 6502 4435 6554
rect 4435 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4261 6500 4317 6502
rect 4341 6500 4397 6502
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 3601 4922 3657 4924
rect 3681 4922 3737 4924
rect 3761 4922 3817 4924
rect 3841 4922 3897 4924
rect 3601 4870 3647 4922
rect 3647 4870 3657 4922
rect 3681 4870 3711 4922
rect 3711 4870 3723 4922
rect 3723 4870 3737 4922
rect 3761 4870 3775 4922
rect 3775 4870 3787 4922
rect 3787 4870 3817 4922
rect 3841 4870 3851 4922
rect 3851 4870 3897 4922
rect 3601 4868 3657 4870
rect 3681 4868 3737 4870
rect 3761 4868 3817 4870
rect 3841 4868 3897 4870
rect 3601 3834 3657 3836
rect 3681 3834 3737 3836
rect 3761 3834 3817 3836
rect 3841 3834 3897 3836
rect 3601 3782 3647 3834
rect 3647 3782 3657 3834
rect 3681 3782 3711 3834
rect 3711 3782 3723 3834
rect 3723 3782 3737 3834
rect 3761 3782 3775 3834
rect 3775 3782 3787 3834
rect 3787 3782 3817 3834
rect 3841 3782 3851 3834
rect 3851 3782 3897 3834
rect 3601 3780 3657 3782
rect 3681 3780 3737 3782
rect 3761 3780 3817 3782
rect 3841 3780 3897 3782
rect 4261 5466 4317 5468
rect 4341 5466 4397 5468
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4261 5414 4307 5466
rect 4307 5414 4317 5466
rect 4341 5414 4371 5466
rect 4371 5414 4383 5466
rect 4383 5414 4397 5466
rect 4421 5414 4435 5466
rect 4435 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4261 5412 4317 5414
rect 4341 5412 4397 5414
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4261 4378 4317 4380
rect 4341 4378 4397 4380
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4261 4326 4307 4378
rect 4307 4326 4317 4378
rect 4341 4326 4371 4378
rect 4371 4326 4383 4378
rect 4383 4326 4397 4378
rect 4421 4326 4435 4378
rect 4435 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4261 4324 4317 4326
rect 4341 4324 4397 4326
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4261 3290 4317 3292
rect 4341 3290 4397 3292
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4261 3238 4307 3290
rect 4307 3238 4317 3290
rect 4341 3238 4371 3290
rect 4371 3238 4383 3290
rect 4383 3238 4397 3290
rect 4421 3238 4435 3290
rect 4435 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4261 3236 4317 3238
rect 4341 3236 4397 3238
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 8891 13626 8947 13628
rect 8971 13626 9027 13628
rect 9051 13626 9107 13628
rect 9131 13626 9187 13628
rect 8891 13574 8937 13626
rect 8937 13574 8947 13626
rect 8971 13574 9001 13626
rect 9001 13574 9013 13626
rect 9013 13574 9027 13626
rect 9051 13574 9065 13626
rect 9065 13574 9077 13626
rect 9077 13574 9107 13626
rect 9131 13574 9141 13626
rect 9141 13574 9187 13626
rect 8891 13572 8947 13574
rect 8971 13572 9027 13574
rect 9051 13572 9107 13574
rect 9131 13572 9187 13574
rect 9551 14170 9607 14172
rect 9631 14170 9687 14172
rect 9711 14170 9767 14172
rect 9791 14170 9847 14172
rect 9551 14118 9597 14170
rect 9597 14118 9607 14170
rect 9631 14118 9661 14170
rect 9661 14118 9673 14170
rect 9673 14118 9687 14170
rect 9711 14118 9725 14170
rect 9725 14118 9737 14170
rect 9737 14118 9767 14170
rect 9791 14118 9801 14170
rect 9801 14118 9847 14170
rect 9551 14116 9607 14118
rect 9631 14116 9687 14118
rect 9711 14116 9767 14118
rect 9791 14116 9847 14118
rect 9551 13082 9607 13084
rect 9631 13082 9687 13084
rect 9711 13082 9767 13084
rect 9791 13082 9847 13084
rect 9551 13030 9597 13082
rect 9597 13030 9607 13082
rect 9631 13030 9661 13082
rect 9661 13030 9673 13082
rect 9673 13030 9687 13082
rect 9711 13030 9725 13082
rect 9725 13030 9737 13082
rect 9737 13030 9767 13082
rect 9791 13030 9801 13082
rect 9801 13030 9847 13082
rect 9551 13028 9607 13030
rect 9631 13028 9687 13030
rect 9711 13028 9767 13030
rect 9791 13028 9847 13030
rect 8891 12538 8947 12540
rect 8971 12538 9027 12540
rect 9051 12538 9107 12540
rect 9131 12538 9187 12540
rect 8891 12486 8937 12538
rect 8937 12486 8947 12538
rect 8971 12486 9001 12538
rect 9001 12486 9013 12538
rect 9013 12486 9027 12538
rect 9051 12486 9065 12538
rect 9065 12486 9077 12538
rect 9077 12486 9107 12538
rect 9131 12486 9141 12538
rect 9141 12486 9187 12538
rect 8891 12484 8947 12486
rect 8971 12484 9027 12486
rect 9051 12484 9107 12486
rect 9131 12484 9187 12486
rect 9551 11994 9607 11996
rect 9631 11994 9687 11996
rect 9711 11994 9767 11996
rect 9791 11994 9847 11996
rect 9551 11942 9597 11994
rect 9597 11942 9607 11994
rect 9631 11942 9661 11994
rect 9661 11942 9673 11994
rect 9673 11942 9687 11994
rect 9711 11942 9725 11994
rect 9725 11942 9737 11994
rect 9737 11942 9767 11994
rect 9791 11942 9801 11994
rect 9801 11942 9847 11994
rect 9551 11940 9607 11942
rect 9631 11940 9687 11942
rect 9711 11940 9767 11942
rect 9791 11940 9847 11942
rect 8891 11450 8947 11452
rect 8971 11450 9027 11452
rect 9051 11450 9107 11452
rect 9131 11450 9187 11452
rect 8891 11398 8937 11450
rect 8937 11398 8947 11450
rect 8971 11398 9001 11450
rect 9001 11398 9013 11450
rect 9013 11398 9027 11450
rect 9051 11398 9065 11450
rect 9065 11398 9077 11450
rect 9077 11398 9107 11450
rect 9131 11398 9141 11450
rect 9141 11398 9187 11450
rect 8891 11396 8947 11398
rect 8971 11396 9027 11398
rect 9051 11396 9107 11398
rect 9131 11396 9187 11398
rect 9551 10906 9607 10908
rect 9631 10906 9687 10908
rect 9711 10906 9767 10908
rect 9791 10906 9847 10908
rect 9551 10854 9597 10906
rect 9597 10854 9607 10906
rect 9631 10854 9661 10906
rect 9661 10854 9673 10906
rect 9673 10854 9687 10906
rect 9711 10854 9725 10906
rect 9725 10854 9737 10906
rect 9737 10854 9767 10906
rect 9791 10854 9801 10906
rect 9801 10854 9847 10906
rect 9551 10852 9607 10854
rect 9631 10852 9687 10854
rect 9711 10852 9767 10854
rect 9791 10852 9847 10854
rect 8891 10362 8947 10364
rect 8971 10362 9027 10364
rect 9051 10362 9107 10364
rect 9131 10362 9187 10364
rect 8891 10310 8937 10362
rect 8937 10310 8947 10362
rect 8971 10310 9001 10362
rect 9001 10310 9013 10362
rect 9013 10310 9027 10362
rect 9051 10310 9065 10362
rect 9065 10310 9077 10362
rect 9077 10310 9107 10362
rect 9131 10310 9141 10362
rect 9141 10310 9187 10362
rect 8891 10308 8947 10310
rect 8971 10308 9027 10310
rect 9051 10308 9107 10310
rect 9131 10308 9187 10310
rect 9551 9818 9607 9820
rect 9631 9818 9687 9820
rect 9711 9818 9767 9820
rect 9791 9818 9847 9820
rect 9551 9766 9597 9818
rect 9597 9766 9607 9818
rect 9631 9766 9661 9818
rect 9661 9766 9673 9818
rect 9673 9766 9687 9818
rect 9711 9766 9725 9818
rect 9725 9766 9737 9818
rect 9737 9766 9767 9818
rect 9791 9766 9801 9818
rect 9801 9766 9847 9818
rect 9551 9764 9607 9766
rect 9631 9764 9687 9766
rect 9711 9764 9767 9766
rect 9791 9764 9847 9766
rect 8891 9274 8947 9276
rect 8971 9274 9027 9276
rect 9051 9274 9107 9276
rect 9131 9274 9187 9276
rect 8891 9222 8937 9274
rect 8937 9222 8947 9274
rect 8971 9222 9001 9274
rect 9001 9222 9013 9274
rect 9013 9222 9027 9274
rect 9051 9222 9065 9274
rect 9065 9222 9077 9274
rect 9077 9222 9107 9274
rect 9131 9222 9141 9274
rect 9141 9222 9187 9274
rect 8891 9220 8947 9222
rect 8971 9220 9027 9222
rect 9051 9220 9107 9222
rect 9131 9220 9187 9222
rect 8891 8186 8947 8188
rect 8971 8186 9027 8188
rect 9051 8186 9107 8188
rect 9131 8186 9187 8188
rect 8891 8134 8937 8186
rect 8937 8134 8947 8186
rect 8971 8134 9001 8186
rect 9001 8134 9013 8186
rect 9013 8134 9027 8186
rect 9051 8134 9065 8186
rect 9065 8134 9077 8186
rect 9077 8134 9107 8186
rect 9131 8134 9141 8186
rect 9141 8134 9187 8186
rect 8891 8132 8947 8134
rect 8971 8132 9027 8134
rect 9051 8132 9107 8134
rect 9131 8132 9187 8134
rect 9551 8730 9607 8732
rect 9631 8730 9687 8732
rect 9711 8730 9767 8732
rect 9791 8730 9847 8732
rect 9551 8678 9597 8730
rect 9597 8678 9607 8730
rect 9631 8678 9661 8730
rect 9661 8678 9673 8730
rect 9673 8678 9687 8730
rect 9711 8678 9725 8730
rect 9725 8678 9737 8730
rect 9737 8678 9767 8730
rect 9791 8678 9801 8730
rect 9801 8678 9847 8730
rect 9551 8676 9607 8678
rect 9631 8676 9687 8678
rect 9711 8676 9767 8678
rect 9791 8676 9847 8678
rect 9862 8508 9864 8528
rect 9864 8508 9916 8528
rect 9916 8508 9918 8528
rect 9862 8472 9918 8508
rect 8891 7098 8947 7100
rect 8971 7098 9027 7100
rect 9051 7098 9107 7100
rect 9131 7098 9187 7100
rect 8891 7046 8937 7098
rect 8937 7046 8947 7098
rect 8971 7046 9001 7098
rect 9001 7046 9013 7098
rect 9013 7046 9027 7098
rect 9051 7046 9065 7098
rect 9065 7046 9077 7098
rect 9077 7046 9107 7098
rect 9131 7046 9141 7098
rect 9141 7046 9187 7098
rect 8891 7044 8947 7046
rect 8971 7044 9027 7046
rect 9051 7044 9107 7046
rect 9131 7044 9187 7046
rect 10230 8472 10286 8528
rect 9551 7642 9607 7644
rect 9631 7642 9687 7644
rect 9711 7642 9767 7644
rect 9791 7642 9847 7644
rect 9551 7590 9597 7642
rect 9597 7590 9607 7642
rect 9631 7590 9661 7642
rect 9661 7590 9673 7642
rect 9673 7590 9687 7642
rect 9711 7590 9725 7642
rect 9725 7590 9737 7642
rect 9737 7590 9767 7642
rect 9791 7590 9801 7642
rect 9801 7590 9847 7642
rect 9551 7588 9607 7590
rect 9631 7588 9687 7590
rect 9711 7588 9767 7590
rect 9791 7588 9847 7590
rect 8891 6010 8947 6012
rect 8971 6010 9027 6012
rect 9051 6010 9107 6012
rect 9131 6010 9187 6012
rect 8891 5958 8937 6010
rect 8937 5958 8947 6010
rect 8971 5958 9001 6010
rect 9001 5958 9013 6010
rect 9013 5958 9027 6010
rect 9051 5958 9065 6010
rect 9065 5958 9077 6010
rect 9077 5958 9107 6010
rect 9131 5958 9141 6010
rect 9141 5958 9187 6010
rect 8891 5956 8947 5958
rect 8971 5956 9027 5958
rect 9051 5956 9107 5958
rect 9131 5956 9187 5958
rect 9551 6554 9607 6556
rect 9631 6554 9687 6556
rect 9711 6554 9767 6556
rect 9791 6554 9847 6556
rect 9551 6502 9597 6554
rect 9597 6502 9607 6554
rect 9631 6502 9661 6554
rect 9661 6502 9673 6554
rect 9673 6502 9687 6554
rect 9711 6502 9725 6554
rect 9725 6502 9737 6554
rect 9737 6502 9767 6554
rect 9791 6502 9801 6554
rect 9801 6502 9847 6554
rect 9551 6500 9607 6502
rect 9631 6500 9687 6502
rect 9711 6500 9767 6502
rect 9791 6500 9847 6502
rect 8891 4922 8947 4924
rect 8971 4922 9027 4924
rect 9051 4922 9107 4924
rect 9131 4922 9187 4924
rect 8891 4870 8937 4922
rect 8937 4870 8947 4922
rect 8971 4870 9001 4922
rect 9001 4870 9013 4922
rect 9013 4870 9027 4922
rect 9051 4870 9065 4922
rect 9065 4870 9077 4922
rect 9077 4870 9107 4922
rect 9131 4870 9141 4922
rect 9141 4870 9187 4922
rect 8891 4868 8947 4870
rect 8971 4868 9027 4870
rect 9051 4868 9107 4870
rect 9131 4868 9187 4870
rect 9678 5636 9734 5672
rect 9678 5616 9680 5636
rect 9680 5616 9732 5636
rect 9732 5616 9734 5636
rect 9551 5466 9607 5468
rect 9631 5466 9687 5468
rect 9711 5466 9767 5468
rect 9791 5466 9847 5468
rect 9551 5414 9597 5466
rect 9597 5414 9607 5466
rect 9631 5414 9661 5466
rect 9661 5414 9673 5466
rect 9673 5414 9687 5466
rect 9711 5414 9725 5466
rect 9725 5414 9737 5466
rect 9737 5414 9767 5466
rect 9791 5414 9801 5466
rect 9801 5414 9847 5466
rect 9551 5412 9607 5414
rect 9631 5412 9687 5414
rect 9711 5412 9767 5414
rect 9791 5412 9847 5414
rect 9551 4378 9607 4380
rect 9631 4378 9687 4380
rect 9711 4378 9767 4380
rect 9791 4378 9847 4380
rect 9551 4326 9597 4378
rect 9597 4326 9607 4378
rect 9631 4326 9661 4378
rect 9661 4326 9673 4378
rect 9673 4326 9687 4378
rect 9711 4326 9725 4378
rect 9725 4326 9737 4378
rect 9737 4326 9767 4378
rect 9791 4326 9801 4378
rect 9801 4326 9847 4378
rect 9551 4324 9607 4326
rect 9631 4324 9687 4326
rect 9711 4324 9767 4326
rect 9791 4324 9847 4326
rect 9770 4156 9772 4176
rect 9772 4156 9824 4176
rect 9824 4156 9826 4176
rect 8891 3834 8947 3836
rect 8971 3834 9027 3836
rect 9051 3834 9107 3836
rect 9131 3834 9187 3836
rect 8891 3782 8937 3834
rect 8937 3782 8947 3834
rect 8971 3782 9001 3834
rect 9001 3782 9013 3834
rect 9013 3782 9027 3834
rect 9051 3782 9065 3834
rect 9065 3782 9077 3834
rect 9077 3782 9107 3834
rect 9131 3782 9141 3834
rect 9141 3782 9187 3834
rect 8891 3780 8947 3782
rect 8971 3780 9027 3782
rect 9051 3780 9107 3782
rect 9131 3780 9187 3782
rect 9770 4120 9826 4156
rect 11886 15544 11942 15600
rect 14181 22330 14237 22332
rect 14261 22330 14317 22332
rect 14341 22330 14397 22332
rect 14421 22330 14477 22332
rect 14181 22278 14227 22330
rect 14227 22278 14237 22330
rect 14261 22278 14291 22330
rect 14291 22278 14303 22330
rect 14303 22278 14317 22330
rect 14341 22278 14355 22330
rect 14355 22278 14367 22330
rect 14367 22278 14397 22330
rect 14421 22278 14431 22330
rect 14431 22278 14477 22330
rect 14181 22276 14237 22278
rect 14261 22276 14317 22278
rect 14341 22276 14397 22278
rect 14421 22276 14477 22278
rect 14841 21786 14897 21788
rect 14921 21786 14977 21788
rect 15001 21786 15057 21788
rect 15081 21786 15137 21788
rect 14841 21734 14887 21786
rect 14887 21734 14897 21786
rect 14921 21734 14951 21786
rect 14951 21734 14963 21786
rect 14963 21734 14977 21786
rect 15001 21734 15015 21786
rect 15015 21734 15027 21786
rect 15027 21734 15057 21786
rect 15081 21734 15091 21786
rect 15091 21734 15137 21786
rect 14841 21732 14897 21734
rect 14921 21732 14977 21734
rect 15001 21732 15057 21734
rect 15081 21732 15137 21734
rect 14181 21242 14237 21244
rect 14261 21242 14317 21244
rect 14341 21242 14397 21244
rect 14421 21242 14477 21244
rect 14181 21190 14227 21242
rect 14227 21190 14237 21242
rect 14261 21190 14291 21242
rect 14291 21190 14303 21242
rect 14303 21190 14317 21242
rect 14341 21190 14355 21242
rect 14355 21190 14367 21242
rect 14367 21190 14397 21242
rect 14421 21190 14431 21242
rect 14431 21190 14477 21242
rect 14181 21188 14237 21190
rect 14261 21188 14317 21190
rect 14341 21188 14397 21190
rect 14421 21188 14477 21190
rect 14841 20698 14897 20700
rect 14921 20698 14977 20700
rect 15001 20698 15057 20700
rect 15081 20698 15137 20700
rect 14841 20646 14887 20698
rect 14887 20646 14897 20698
rect 14921 20646 14951 20698
rect 14951 20646 14963 20698
rect 14963 20646 14977 20698
rect 15001 20646 15015 20698
rect 15015 20646 15027 20698
rect 15027 20646 15057 20698
rect 15081 20646 15091 20698
rect 15091 20646 15137 20698
rect 14841 20644 14897 20646
rect 14921 20644 14977 20646
rect 15001 20644 15057 20646
rect 15081 20644 15137 20646
rect 16302 21292 16304 21312
rect 16304 21292 16356 21312
rect 16356 21292 16358 21312
rect 16302 21256 16358 21292
rect 14181 20154 14237 20156
rect 14261 20154 14317 20156
rect 14341 20154 14397 20156
rect 14421 20154 14477 20156
rect 14181 20102 14227 20154
rect 14227 20102 14237 20154
rect 14261 20102 14291 20154
rect 14291 20102 14303 20154
rect 14303 20102 14317 20154
rect 14341 20102 14355 20154
rect 14355 20102 14367 20154
rect 14367 20102 14397 20154
rect 14421 20102 14431 20154
rect 14431 20102 14477 20154
rect 14181 20100 14237 20102
rect 14261 20100 14317 20102
rect 14341 20100 14397 20102
rect 14421 20100 14477 20102
rect 14841 19610 14897 19612
rect 14921 19610 14977 19612
rect 15001 19610 15057 19612
rect 15081 19610 15137 19612
rect 14841 19558 14887 19610
rect 14887 19558 14897 19610
rect 14921 19558 14951 19610
rect 14951 19558 14963 19610
rect 14963 19558 14977 19610
rect 15001 19558 15015 19610
rect 15015 19558 15027 19610
rect 15027 19558 15057 19610
rect 15081 19558 15091 19610
rect 15091 19558 15137 19610
rect 14841 19556 14897 19558
rect 14921 19556 14977 19558
rect 15001 19556 15057 19558
rect 15081 19556 15137 19558
rect 14181 19066 14237 19068
rect 14261 19066 14317 19068
rect 14341 19066 14397 19068
rect 14421 19066 14477 19068
rect 14181 19014 14227 19066
rect 14227 19014 14237 19066
rect 14261 19014 14291 19066
rect 14291 19014 14303 19066
rect 14303 19014 14317 19066
rect 14341 19014 14355 19066
rect 14355 19014 14367 19066
rect 14367 19014 14397 19066
rect 14421 19014 14431 19066
rect 14431 19014 14477 19066
rect 14181 19012 14237 19014
rect 14261 19012 14317 19014
rect 14341 19012 14397 19014
rect 14421 19012 14477 19014
rect 14002 18164 14004 18184
rect 14004 18164 14056 18184
rect 14056 18164 14058 18184
rect 14002 18128 14058 18164
rect 14841 18522 14897 18524
rect 14921 18522 14977 18524
rect 15001 18522 15057 18524
rect 15081 18522 15137 18524
rect 14841 18470 14887 18522
rect 14887 18470 14897 18522
rect 14921 18470 14951 18522
rect 14951 18470 14963 18522
rect 14963 18470 14977 18522
rect 15001 18470 15015 18522
rect 15015 18470 15027 18522
rect 15027 18470 15057 18522
rect 15081 18470 15091 18522
rect 15091 18470 15137 18522
rect 14841 18468 14897 18470
rect 14921 18468 14977 18470
rect 15001 18468 15057 18470
rect 15081 18468 15137 18470
rect 14181 17978 14237 17980
rect 14261 17978 14317 17980
rect 14341 17978 14397 17980
rect 14421 17978 14477 17980
rect 14181 17926 14227 17978
rect 14227 17926 14237 17978
rect 14261 17926 14291 17978
rect 14291 17926 14303 17978
rect 14303 17926 14317 17978
rect 14341 17926 14355 17978
rect 14355 17926 14367 17978
rect 14367 17926 14397 17978
rect 14421 17926 14431 17978
rect 14431 17926 14477 17978
rect 14181 17924 14237 17926
rect 14261 17924 14317 17926
rect 14341 17924 14397 17926
rect 14421 17924 14477 17926
rect 14841 17434 14897 17436
rect 14921 17434 14977 17436
rect 15001 17434 15057 17436
rect 15081 17434 15137 17436
rect 14841 17382 14887 17434
rect 14887 17382 14897 17434
rect 14921 17382 14951 17434
rect 14951 17382 14963 17434
rect 14963 17382 14977 17434
rect 15001 17382 15015 17434
rect 15015 17382 15027 17434
rect 15027 17382 15057 17434
rect 15081 17382 15091 17434
rect 15091 17382 15137 17434
rect 14841 17380 14897 17382
rect 14921 17380 14977 17382
rect 15001 17380 15057 17382
rect 15081 17380 15137 17382
rect 14181 16890 14237 16892
rect 14261 16890 14317 16892
rect 14341 16890 14397 16892
rect 14421 16890 14477 16892
rect 14181 16838 14227 16890
rect 14227 16838 14237 16890
rect 14261 16838 14291 16890
rect 14291 16838 14303 16890
rect 14303 16838 14317 16890
rect 14341 16838 14355 16890
rect 14355 16838 14367 16890
rect 14367 16838 14397 16890
rect 14421 16838 14431 16890
rect 14431 16838 14477 16890
rect 14181 16836 14237 16838
rect 14261 16836 14317 16838
rect 14341 16836 14397 16838
rect 14421 16836 14477 16838
rect 14181 15802 14237 15804
rect 14261 15802 14317 15804
rect 14341 15802 14397 15804
rect 14421 15802 14477 15804
rect 14181 15750 14227 15802
rect 14227 15750 14237 15802
rect 14261 15750 14291 15802
rect 14291 15750 14303 15802
rect 14303 15750 14317 15802
rect 14341 15750 14355 15802
rect 14355 15750 14367 15802
rect 14367 15750 14397 15802
rect 14421 15750 14431 15802
rect 14431 15750 14477 15802
rect 14181 15748 14237 15750
rect 14261 15748 14317 15750
rect 14341 15748 14397 15750
rect 14421 15748 14477 15750
rect 14841 16346 14897 16348
rect 14921 16346 14977 16348
rect 15001 16346 15057 16348
rect 15081 16346 15137 16348
rect 14841 16294 14887 16346
rect 14887 16294 14897 16346
rect 14921 16294 14951 16346
rect 14951 16294 14963 16346
rect 14963 16294 14977 16346
rect 15001 16294 15015 16346
rect 15015 16294 15027 16346
rect 15027 16294 15057 16346
rect 15081 16294 15091 16346
rect 15091 16294 15137 16346
rect 14841 16292 14897 16294
rect 14921 16292 14977 16294
rect 15001 16292 15057 16294
rect 15081 16292 15137 16294
rect 15290 15544 15346 15600
rect 14841 15258 14897 15260
rect 14921 15258 14977 15260
rect 15001 15258 15057 15260
rect 15081 15258 15137 15260
rect 14841 15206 14887 15258
rect 14887 15206 14897 15258
rect 14921 15206 14951 15258
rect 14951 15206 14963 15258
rect 14963 15206 14977 15258
rect 15001 15206 15015 15258
rect 15015 15206 15027 15258
rect 15027 15206 15057 15258
rect 15081 15206 15091 15258
rect 15091 15206 15137 15258
rect 14841 15204 14897 15206
rect 14921 15204 14977 15206
rect 15001 15204 15057 15206
rect 15081 15204 15137 15206
rect 14181 14714 14237 14716
rect 14261 14714 14317 14716
rect 14341 14714 14397 14716
rect 14421 14714 14477 14716
rect 14181 14662 14227 14714
rect 14227 14662 14237 14714
rect 14261 14662 14291 14714
rect 14291 14662 14303 14714
rect 14303 14662 14317 14714
rect 14341 14662 14355 14714
rect 14355 14662 14367 14714
rect 14367 14662 14397 14714
rect 14421 14662 14431 14714
rect 14431 14662 14477 14714
rect 14181 14660 14237 14662
rect 14261 14660 14317 14662
rect 14341 14660 14397 14662
rect 14421 14660 14477 14662
rect 14841 14170 14897 14172
rect 14921 14170 14977 14172
rect 15001 14170 15057 14172
rect 15081 14170 15137 14172
rect 14841 14118 14887 14170
rect 14887 14118 14897 14170
rect 14921 14118 14951 14170
rect 14951 14118 14963 14170
rect 14963 14118 14977 14170
rect 15001 14118 15015 14170
rect 15015 14118 15027 14170
rect 15027 14118 15057 14170
rect 15081 14118 15091 14170
rect 15091 14118 15137 14170
rect 14841 14116 14897 14118
rect 14921 14116 14977 14118
rect 15001 14116 15057 14118
rect 15081 14116 15137 14118
rect 15566 18128 15622 18184
rect 16946 21256 17002 21312
rect 16578 19352 16634 19408
rect 19471 22330 19527 22332
rect 19551 22330 19607 22332
rect 19631 22330 19687 22332
rect 19711 22330 19767 22332
rect 19471 22278 19517 22330
rect 19517 22278 19527 22330
rect 19551 22278 19581 22330
rect 19581 22278 19593 22330
rect 19593 22278 19607 22330
rect 19631 22278 19645 22330
rect 19645 22278 19657 22330
rect 19657 22278 19687 22330
rect 19711 22278 19721 22330
rect 19721 22278 19767 22330
rect 19471 22276 19527 22278
rect 19551 22276 19607 22278
rect 19631 22276 19687 22278
rect 19711 22276 19767 22278
rect 20131 21786 20187 21788
rect 20211 21786 20267 21788
rect 20291 21786 20347 21788
rect 20371 21786 20427 21788
rect 20131 21734 20177 21786
rect 20177 21734 20187 21786
rect 20211 21734 20241 21786
rect 20241 21734 20253 21786
rect 20253 21734 20267 21786
rect 20291 21734 20305 21786
rect 20305 21734 20317 21786
rect 20317 21734 20347 21786
rect 20371 21734 20381 21786
rect 20381 21734 20427 21786
rect 20131 21732 20187 21734
rect 20211 21732 20267 21734
rect 20291 21732 20347 21734
rect 20371 21732 20427 21734
rect 19471 21242 19527 21244
rect 19551 21242 19607 21244
rect 19631 21242 19687 21244
rect 19711 21242 19767 21244
rect 19471 21190 19517 21242
rect 19517 21190 19527 21242
rect 19551 21190 19581 21242
rect 19581 21190 19593 21242
rect 19593 21190 19607 21242
rect 19631 21190 19645 21242
rect 19645 21190 19657 21242
rect 19657 21190 19687 21242
rect 19711 21190 19721 21242
rect 19721 21190 19767 21242
rect 19471 21188 19527 21190
rect 19551 21188 19607 21190
rect 19631 21188 19687 21190
rect 19711 21188 19767 21190
rect 20131 20698 20187 20700
rect 20211 20698 20267 20700
rect 20291 20698 20347 20700
rect 20371 20698 20427 20700
rect 20131 20646 20177 20698
rect 20177 20646 20187 20698
rect 20211 20646 20241 20698
rect 20241 20646 20253 20698
rect 20253 20646 20267 20698
rect 20291 20646 20305 20698
rect 20305 20646 20317 20698
rect 20317 20646 20347 20698
rect 20371 20646 20381 20698
rect 20381 20646 20427 20698
rect 20131 20644 20187 20646
rect 20211 20644 20267 20646
rect 20291 20644 20347 20646
rect 20371 20644 20427 20646
rect 22190 21120 22246 21176
rect 19471 20154 19527 20156
rect 19551 20154 19607 20156
rect 19631 20154 19687 20156
rect 19711 20154 19767 20156
rect 19471 20102 19517 20154
rect 19517 20102 19527 20154
rect 19551 20102 19581 20154
rect 19581 20102 19593 20154
rect 19593 20102 19607 20154
rect 19631 20102 19645 20154
rect 19645 20102 19657 20154
rect 19657 20102 19687 20154
rect 19711 20102 19721 20154
rect 19721 20102 19767 20154
rect 19471 20100 19527 20102
rect 19551 20100 19607 20102
rect 19631 20100 19687 20102
rect 19711 20100 19767 20102
rect 20131 19610 20187 19612
rect 20211 19610 20267 19612
rect 20291 19610 20347 19612
rect 20371 19610 20427 19612
rect 20131 19558 20177 19610
rect 20177 19558 20187 19610
rect 20211 19558 20241 19610
rect 20241 19558 20253 19610
rect 20253 19558 20267 19610
rect 20291 19558 20305 19610
rect 20305 19558 20317 19610
rect 20317 19558 20347 19610
rect 20371 19558 20381 19610
rect 20381 19558 20427 19610
rect 20131 19556 20187 19558
rect 20211 19556 20267 19558
rect 20291 19556 20347 19558
rect 20371 19556 20427 19558
rect 19471 19066 19527 19068
rect 19551 19066 19607 19068
rect 19631 19066 19687 19068
rect 19711 19066 19767 19068
rect 19471 19014 19517 19066
rect 19517 19014 19527 19066
rect 19551 19014 19581 19066
rect 19581 19014 19593 19066
rect 19593 19014 19607 19066
rect 19631 19014 19645 19066
rect 19645 19014 19657 19066
rect 19657 19014 19687 19066
rect 19711 19014 19721 19066
rect 19721 19014 19767 19066
rect 19471 19012 19527 19014
rect 19551 19012 19607 19014
rect 19631 19012 19687 19014
rect 19711 19012 19767 19014
rect 20131 18522 20187 18524
rect 20211 18522 20267 18524
rect 20291 18522 20347 18524
rect 20371 18522 20427 18524
rect 20131 18470 20177 18522
rect 20177 18470 20187 18522
rect 20211 18470 20241 18522
rect 20241 18470 20253 18522
rect 20253 18470 20267 18522
rect 20291 18470 20305 18522
rect 20305 18470 20317 18522
rect 20317 18470 20347 18522
rect 20371 18470 20381 18522
rect 20381 18470 20427 18522
rect 20131 18468 20187 18470
rect 20211 18468 20267 18470
rect 20291 18468 20347 18470
rect 20371 18468 20427 18470
rect 19471 17978 19527 17980
rect 19551 17978 19607 17980
rect 19631 17978 19687 17980
rect 19711 17978 19767 17980
rect 19471 17926 19517 17978
rect 19517 17926 19527 17978
rect 19551 17926 19581 17978
rect 19581 17926 19593 17978
rect 19593 17926 19607 17978
rect 19631 17926 19645 17978
rect 19645 17926 19657 17978
rect 19657 17926 19687 17978
rect 19711 17926 19721 17978
rect 19721 17926 19767 17978
rect 19471 17924 19527 17926
rect 19551 17924 19607 17926
rect 19631 17924 19687 17926
rect 19711 17924 19767 17926
rect 19471 16890 19527 16892
rect 19551 16890 19607 16892
rect 19631 16890 19687 16892
rect 19711 16890 19767 16892
rect 19471 16838 19517 16890
rect 19517 16838 19527 16890
rect 19551 16838 19581 16890
rect 19581 16838 19593 16890
rect 19593 16838 19607 16890
rect 19631 16838 19645 16890
rect 19645 16838 19657 16890
rect 19657 16838 19687 16890
rect 19711 16838 19721 16890
rect 19721 16838 19767 16890
rect 19471 16836 19527 16838
rect 19551 16836 19607 16838
rect 19631 16836 19687 16838
rect 19711 16836 19767 16838
rect 20131 17434 20187 17436
rect 20211 17434 20267 17436
rect 20291 17434 20347 17436
rect 20371 17434 20427 17436
rect 20131 17382 20177 17434
rect 20177 17382 20187 17434
rect 20211 17382 20241 17434
rect 20241 17382 20253 17434
rect 20253 17382 20267 17434
rect 20291 17382 20305 17434
rect 20305 17382 20317 17434
rect 20317 17382 20347 17434
rect 20371 17382 20381 17434
rect 20381 17382 20427 17434
rect 20131 17380 20187 17382
rect 20211 17380 20267 17382
rect 20291 17380 20347 17382
rect 20371 17380 20427 17382
rect 14181 13626 14237 13628
rect 14261 13626 14317 13628
rect 14341 13626 14397 13628
rect 14421 13626 14477 13628
rect 14181 13574 14227 13626
rect 14227 13574 14237 13626
rect 14261 13574 14291 13626
rect 14291 13574 14303 13626
rect 14303 13574 14317 13626
rect 14341 13574 14355 13626
rect 14355 13574 14367 13626
rect 14367 13574 14397 13626
rect 14421 13574 14431 13626
rect 14431 13574 14477 13626
rect 14181 13572 14237 13574
rect 14261 13572 14317 13574
rect 14341 13572 14397 13574
rect 14421 13572 14477 13574
rect 14841 13082 14897 13084
rect 14921 13082 14977 13084
rect 15001 13082 15057 13084
rect 15081 13082 15137 13084
rect 14841 13030 14887 13082
rect 14887 13030 14897 13082
rect 14921 13030 14951 13082
rect 14951 13030 14963 13082
rect 14963 13030 14977 13082
rect 15001 13030 15015 13082
rect 15015 13030 15027 13082
rect 15027 13030 15057 13082
rect 15081 13030 15091 13082
rect 15091 13030 15137 13082
rect 14841 13028 14897 13030
rect 14921 13028 14977 13030
rect 15001 13028 15057 13030
rect 15081 13028 15137 13030
rect 14181 12538 14237 12540
rect 14261 12538 14317 12540
rect 14341 12538 14397 12540
rect 14421 12538 14477 12540
rect 14181 12486 14227 12538
rect 14227 12486 14237 12538
rect 14261 12486 14291 12538
rect 14291 12486 14303 12538
rect 14303 12486 14317 12538
rect 14341 12486 14355 12538
rect 14355 12486 14367 12538
rect 14367 12486 14397 12538
rect 14421 12486 14431 12538
rect 14431 12486 14477 12538
rect 14181 12484 14237 12486
rect 14261 12484 14317 12486
rect 14341 12484 14397 12486
rect 14421 12484 14477 12486
rect 14181 11450 14237 11452
rect 14261 11450 14317 11452
rect 14341 11450 14397 11452
rect 14421 11450 14477 11452
rect 14181 11398 14227 11450
rect 14227 11398 14237 11450
rect 14261 11398 14291 11450
rect 14291 11398 14303 11450
rect 14303 11398 14317 11450
rect 14341 11398 14355 11450
rect 14355 11398 14367 11450
rect 14367 11398 14397 11450
rect 14421 11398 14431 11450
rect 14431 11398 14477 11450
rect 14181 11396 14237 11398
rect 14261 11396 14317 11398
rect 14341 11396 14397 11398
rect 14421 11396 14477 11398
rect 14181 10362 14237 10364
rect 14261 10362 14317 10364
rect 14341 10362 14397 10364
rect 14421 10362 14477 10364
rect 14181 10310 14227 10362
rect 14227 10310 14237 10362
rect 14261 10310 14291 10362
rect 14291 10310 14303 10362
rect 14303 10310 14317 10362
rect 14341 10310 14355 10362
rect 14355 10310 14367 10362
rect 14367 10310 14397 10362
rect 14421 10310 14431 10362
rect 14431 10310 14477 10362
rect 14181 10308 14237 10310
rect 14261 10308 14317 10310
rect 14341 10308 14397 10310
rect 14421 10308 14477 10310
rect 11518 8472 11574 8528
rect 14181 9274 14237 9276
rect 14261 9274 14317 9276
rect 14341 9274 14397 9276
rect 14421 9274 14477 9276
rect 14181 9222 14227 9274
rect 14227 9222 14237 9274
rect 14261 9222 14291 9274
rect 14291 9222 14303 9274
rect 14303 9222 14317 9274
rect 14341 9222 14355 9274
rect 14355 9222 14367 9274
rect 14367 9222 14397 9274
rect 14421 9222 14431 9274
rect 14431 9222 14477 9274
rect 14181 9220 14237 9222
rect 14261 9220 14317 9222
rect 14341 9220 14397 9222
rect 14421 9220 14477 9222
rect 11150 5652 11152 5672
rect 11152 5652 11204 5672
rect 11204 5652 11206 5672
rect 11150 5616 11206 5652
rect 9551 3290 9607 3292
rect 9631 3290 9687 3292
rect 9711 3290 9767 3292
rect 9791 3290 9847 3292
rect 9551 3238 9597 3290
rect 9597 3238 9607 3290
rect 9631 3238 9661 3290
rect 9661 3238 9673 3290
rect 9673 3238 9687 3290
rect 9711 3238 9725 3290
rect 9725 3238 9737 3290
rect 9737 3238 9767 3290
rect 9791 3238 9801 3290
rect 9801 3238 9847 3290
rect 9551 3236 9607 3238
rect 9631 3236 9687 3238
rect 9711 3236 9767 3238
rect 9791 3236 9847 3238
rect 14181 8186 14237 8188
rect 14261 8186 14317 8188
rect 14341 8186 14397 8188
rect 14421 8186 14477 8188
rect 14181 8134 14227 8186
rect 14227 8134 14237 8186
rect 14261 8134 14291 8186
rect 14291 8134 14303 8186
rect 14303 8134 14317 8186
rect 14341 8134 14355 8186
rect 14355 8134 14367 8186
rect 14367 8134 14397 8186
rect 14421 8134 14431 8186
rect 14431 8134 14477 8186
rect 14181 8132 14237 8134
rect 14261 8132 14317 8134
rect 14341 8132 14397 8134
rect 14421 8132 14477 8134
rect 14181 7098 14237 7100
rect 14261 7098 14317 7100
rect 14341 7098 14397 7100
rect 14421 7098 14477 7100
rect 14181 7046 14227 7098
rect 14227 7046 14237 7098
rect 14261 7046 14291 7098
rect 14291 7046 14303 7098
rect 14303 7046 14317 7098
rect 14341 7046 14355 7098
rect 14355 7046 14367 7098
rect 14367 7046 14397 7098
rect 14421 7046 14431 7098
rect 14431 7046 14477 7098
rect 14181 7044 14237 7046
rect 14261 7044 14317 7046
rect 14341 7044 14397 7046
rect 14421 7044 14477 7046
rect 14181 6010 14237 6012
rect 14261 6010 14317 6012
rect 14341 6010 14397 6012
rect 14421 6010 14477 6012
rect 14181 5958 14227 6010
rect 14227 5958 14237 6010
rect 14261 5958 14291 6010
rect 14291 5958 14303 6010
rect 14303 5958 14317 6010
rect 14341 5958 14355 6010
rect 14355 5958 14367 6010
rect 14367 5958 14397 6010
rect 14421 5958 14431 6010
rect 14431 5958 14477 6010
rect 14181 5956 14237 5958
rect 14261 5956 14317 5958
rect 14341 5956 14397 5958
rect 14421 5956 14477 5958
rect 14841 11994 14897 11996
rect 14921 11994 14977 11996
rect 15001 11994 15057 11996
rect 15081 11994 15137 11996
rect 14841 11942 14887 11994
rect 14887 11942 14897 11994
rect 14921 11942 14951 11994
rect 14951 11942 14963 11994
rect 14963 11942 14977 11994
rect 15001 11942 15015 11994
rect 15015 11942 15027 11994
rect 15027 11942 15057 11994
rect 15081 11942 15091 11994
rect 15091 11942 15137 11994
rect 14841 11940 14897 11942
rect 14921 11940 14977 11942
rect 15001 11940 15057 11942
rect 15081 11940 15137 11942
rect 19614 15972 19670 16008
rect 19614 15952 19616 15972
rect 19616 15952 19668 15972
rect 19668 15952 19670 15972
rect 19471 15802 19527 15804
rect 19551 15802 19607 15804
rect 19631 15802 19687 15804
rect 19711 15802 19767 15804
rect 19471 15750 19517 15802
rect 19517 15750 19527 15802
rect 19551 15750 19581 15802
rect 19581 15750 19593 15802
rect 19593 15750 19607 15802
rect 19631 15750 19645 15802
rect 19645 15750 19657 15802
rect 19657 15750 19687 15802
rect 19711 15750 19721 15802
rect 19721 15750 19767 15802
rect 19471 15748 19527 15750
rect 19551 15748 19607 15750
rect 19631 15748 19687 15750
rect 19711 15748 19767 15750
rect 19338 15544 19394 15600
rect 14841 10906 14897 10908
rect 14921 10906 14977 10908
rect 15001 10906 15057 10908
rect 15081 10906 15137 10908
rect 14841 10854 14887 10906
rect 14887 10854 14897 10906
rect 14921 10854 14951 10906
rect 14951 10854 14963 10906
rect 14963 10854 14977 10906
rect 15001 10854 15015 10906
rect 15015 10854 15027 10906
rect 15027 10854 15057 10906
rect 15081 10854 15091 10906
rect 15091 10854 15137 10906
rect 14841 10852 14897 10854
rect 14921 10852 14977 10854
rect 15001 10852 15057 10854
rect 15081 10852 15137 10854
rect 14841 9818 14897 9820
rect 14921 9818 14977 9820
rect 15001 9818 15057 9820
rect 15081 9818 15137 9820
rect 14841 9766 14887 9818
rect 14887 9766 14897 9818
rect 14921 9766 14951 9818
rect 14951 9766 14963 9818
rect 14963 9766 14977 9818
rect 15001 9766 15015 9818
rect 15015 9766 15027 9818
rect 15027 9766 15057 9818
rect 15081 9766 15091 9818
rect 15091 9766 15137 9818
rect 14841 9764 14897 9766
rect 14921 9764 14977 9766
rect 15001 9764 15057 9766
rect 15081 9764 15137 9766
rect 14841 8730 14897 8732
rect 14921 8730 14977 8732
rect 15001 8730 15057 8732
rect 15081 8730 15137 8732
rect 14841 8678 14887 8730
rect 14887 8678 14897 8730
rect 14921 8678 14951 8730
rect 14951 8678 14963 8730
rect 14963 8678 14977 8730
rect 15001 8678 15015 8730
rect 15015 8678 15027 8730
rect 15027 8678 15057 8730
rect 15081 8678 15091 8730
rect 15091 8678 15137 8730
rect 14841 8676 14897 8678
rect 14921 8676 14977 8678
rect 15001 8676 15057 8678
rect 15081 8676 15137 8678
rect 14841 7642 14897 7644
rect 14921 7642 14977 7644
rect 15001 7642 15057 7644
rect 15081 7642 15137 7644
rect 14841 7590 14887 7642
rect 14887 7590 14897 7642
rect 14921 7590 14951 7642
rect 14951 7590 14963 7642
rect 14963 7590 14977 7642
rect 15001 7590 15015 7642
rect 15015 7590 15027 7642
rect 15027 7590 15057 7642
rect 15081 7590 15091 7642
rect 15091 7590 15137 7642
rect 14841 7588 14897 7590
rect 14921 7588 14977 7590
rect 15001 7588 15057 7590
rect 15081 7588 15137 7590
rect 20074 16496 20130 16552
rect 20131 16346 20187 16348
rect 20211 16346 20267 16348
rect 20291 16346 20347 16348
rect 20371 16346 20427 16348
rect 20131 16294 20177 16346
rect 20177 16294 20187 16346
rect 20211 16294 20241 16346
rect 20241 16294 20253 16346
rect 20253 16294 20267 16346
rect 20291 16294 20305 16346
rect 20305 16294 20317 16346
rect 20317 16294 20347 16346
rect 20371 16294 20381 16346
rect 20381 16294 20427 16346
rect 20131 16292 20187 16294
rect 20211 16292 20267 16294
rect 20291 16292 20347 16294
rect 20371 16292 20427 16294
rect 19982 16088 20038 16144
rect 20131 15258 20187 15260
rect 20211 15258 20267 15260
rect 20291 15258 20347 15260
rect 20371 15258 20427 15260
rect 20131 15206 20177 15258
rect 20177 15206 20187 15258
rect 20211 15206 20241 15258
rect 20241 15206 20253 15258
rect 20253 15206 20267 15258
rect 20291 15206 20305 15258
rect 20305 15206 20317 15258
rect 20317 15206 20347 15258
rect 20371 15206 20381 15258
rect 20381 15206 20427 15258
rect 20131 15204 20187 15206
rect 20211 15204 20267 15206
rect 20291 15204 20347 15206
rect 20371 15204 20427 15206
rect 19471 14714 19527 14716
rect 19551 14714 19607 14716
rect 19631 14714 19687 14716
rect 19711 14714 19767 14716
rect 19471 14662 19517 14714
rect 19517 14662 19527 14714
rect 19551 14662 19581 14714
rect 19581 14662 19593 14714
rect 19593 14662 19607 14714
rect 19631 14662 19645 14714
rect 19645 14662 19657 14714
rect 19657 14662 19687 14714
rect 19711 14662 19721 14714
rect 19721 14662 19767 14714
rect 19471 14660 19527 14662
rect 19551 14660 19607 14662
rect 19631 14660 19687 14662
rect 19711 14660 19767 14662
rect 19471 13626 19527 13628
rect 19551 13626 19607 13628
rect 19631 13626 19687 13628
rect 19711 13626 19767 13628
rect 19471 13574 19517 13626
rect 19517 13574 19527 13626
rect 19551 13574 19581 13626
rect 19581 13574 19593 13626
rect 19593 13574 19607 13626
rect 19631 13574 19645 13626
rect 19645 13574 19657 13626
rect 19657 13574 19687 13626
rect 19711 13574 19721 13626
rect 19721 13574 19767 13626
rect 19471 13572 19527 13574
rect 19551 13572 19607 13574
rect 19631 13572 19687 13574
rect 19711 13572 19767 13574
rect 19471 12538 19527 12540
rect 19551 12538 19607 12540
rect 19631 12538 19687 12540
rect 19711 12538 19767 12540
rect 19471 12486 19517 12538
rect 19517 12486 19527 12538
rect 19551 12486 19581 12538
rect 19581 12486 19593 12538
rect 19593 12486 19607 12538
rect 19631 12486 19645 12538
rect 19645 12486 19657 12538
rect 19657 12486 19687 12538
rect 19711 12486 19721 12538
rect 19721 12486 19767 12538
rect 19471 12484 19527 12486
rect 19551 12484 19607 12486
rect 19631 12484 19687 12486
rect 19711 12484 19767 12486
rect 20131 14170 20187 14172
rect 20211 14170 20267 14172
rect 20291 14170 20347 14172
rect 20371 14170 20427 14172
rect 20131 14118 20177 14170
rect 20177 14118 20187 14170
rect 20211 14118 20241 14170
rect 20241 14118 20253 14170
rect 20253 14118 20267 14170
rect 20291 14118 20305 14170
rect 20305 14118 20317 14170
rect 20317 14118 20347 14170
rect 20371 14118 20381 14170
rect 20381 14118 20427 14170
rect 20131 14116 20187 14118
rect 20211 14116 20267 14118
rect 20291 14116 20347 14118
rect 20371 14116 20427 14118
rect 20131 13082 20187 13084
rect 20211 13082 20267 13084
rect 20291 13082 20347 13084
rect 20371 13082 20427 13084
rect 20131 13030 20177 13082
rect 20177 13030 20187 13082
rect 20211 13030 20241 13082
rect 20241 13030 20253 13082
rect 20253 13030 20267 13082
rect 20291 13030 20305 13082
rect 20305 13030 20317 13082
rect 20317 13030 20347 13082
rect 20371 13030 20381 13082
rect 20381 13030 20427 13082
rect 20131 13028 20187 13030
rect 20211 13028 20267 13030
rect 20291 13028 20347 13030
rect 20371 13028 20427 13030
rect 19471 11450 19527 11452
rect 19551 11450 19607 11452
rect 19631 11450 19687 11452
rect 19711 11450 19767 11452
rect 19471 11398 19517 11450
rect 19517 11398 19527 11450
rect 19551 11398 19581 11450
rect 19581 11398 19593 11450
rect 19593 11398 19607 11450
rect 19631 11398 19645 11450
rect 19645 11398 19657 11450
rect 19657 11398 19687 11450
rect 19711 11398 19721 11450
rect 19721 11398 19767 11450
rect 19471 11396 19527 11398
rect 19551 11396 19607 11398
rect 19631 11396 19687 11398
rect 19711 11396 19767 11398
rect 19471 10362 19527 10364
rect 19551 10362 19607 10364
rect 19631 10362 19687 10364
rect 19711 10362 19767 10364
rect 19471 10310 19517 10362
rect 19517 10310 19527 10362
rect 19551 10310 19581 10362
rect 19581 10310 19593 10362
rect 19593 10310 19607 10362
rect 19631 10310 19645 10362
rect 19645 10310 19657 10362
rect 19657 10310 19687 10362
rect 19711 10310 19721 10362
rect 19721 10310 19767 10362
rect 19471 10308 19527 10310
rect 19551 10308 19607 10310
rect 19631 10308 19687 10310
rect 19711 10308 19767 10310
rect 14841 6554 14897 6556
rect 14921 6554 14977 6556
rect 15001 6554 15057 6556
rect 15081 6554 15137 6556
rect 14841 6502 14887 6554
rect 14887 6502 14897 6554
rect 14921 6502 14951 6554
rect 14951 6502 14963 6554
rect 14963 6502 14977 6554
rect 15001 6502 15015 6554
rect 15015 6502 15027 6554
rect 15027 6502 15057 6554
rect 15081 6502 15091 6554
rect 15091 6502 15137 6554
rect 14841 6500 14897 6502
rect 14921 6500 14977 6502
rect 15001 6500 15057 6502
rect 15081 6500 15137 6502
rect 14841 5466 14897 5468
rect 14921 5466 14977 5468
rect 15001 5466 15057 5468
rect 15081 5466 15137 5468
rect 14841 5414 14887 5466
rect 14887 5414 14897 5466
rect 14921 5414 14951 5466
rect 14951 5414 14963 5466
rect 14963 5414 14977 5466
rect 15001 5414 15015 5466
rect 15015 5414 15027 5466
rect 15027 5414 15057 5466
rect 15081 5414 15091 5466
rect 15091 5414 15137 5466
rect 14841 5412 14897 5414
rect 14921 5412 14977 5414
rect 15001 5412 15057 5414
rect 15081 5412 15137 5414
rect 14181 4922 14237 4924
rect 14261 4922 14317 4924
rect 14341 4922 14397 4924
rect 14421 4922 14477 4924
rect 14181 4870 14227 4922
rect 14227 4870 14237 4922
rect 14261 4870 14291 4922
rect 14291 4870 14303 4922
rect 14303 4870 14317 4922
rect 14341 4870 14355 4922
rect 14355 4870 14367 4922
rect 14367 4870 14397 4922
rect 14421 4870 14431 4922
rect 14431 4870 14477 4922
rect 14181 4868 14237 4870
rect 14261 4868 14317 4870
rect 14341 4868 14397 4870
rect 14421 4868 14477 4870
rect 12990 4120 13046 4176
rect 14841 4378 14897 4380
rect 14921 4378 14977 4380
rect 15001 4378 15057 4380
rect 15081 4378 15137 4380
rect 14841 4326 14887 4378
rect 14887 4326 14897 4378
rect 14921 4326 14951 4378
rect 14951 4326 14963 4378
rect 14963 4326 14977 4378
rect 15001 4326 15015 4378
rect 15015 4326 15027 4378
rect 15027 4326 15057 4378
rect 15081 4326 15091 4378
rect 15091 4326 15137 4378
rect 14841 4324 14897 4326
rect 14921 4324 14977 4326
rect 15001 4324 15057 4326
rect 15081 4324 15137 4326
rect 19471 9274 19527 9276
rect 19551 9274 19607 9276
rect 19631 9274 19687 9276
rect 19711 9274 19767 9276
rect 19471 9222 19517 9274
rect 19517 9222 19527 9274
rect 19551 9222 19581 9274
rect 19581 9222 19593 9274
rect 19593 9222 19607 9274
rect 19631 9222 19645 9274
rect 19645 9222 19657 9274
rect 19657 9222 19687 9274
rect 19711 9222 19721 9274
rect 19721 9222 19767 9274
rect 19471 9220 19527 9222
rect 19551 9220 19607 9222
rect 19631 9220 19687 9222
rect 19711 9220 19767 9222
rect 20131 11994 20187 11996
rect 20211 11994 20267 11996
rect 20291 11994 20347 11996
rect 20371 11994 20427 11996
rect 20131 11942 20177 11994
rect 20177 11942 20187 11994
rect 20211 11942 20241 11994
rect 20241 11942 20253 11994
rect 20253 11942 20267 11994
rect 20291 11942 20305 11994
rect 20305 11942 20317 11994
rect 20317 11942 20347 11994
rect 20371 11942 20381 11994
rect 20381 11942 20427 11994
rect 20131 11940 20187 11942
rect 20211 11940 20267 11942
rect 20291 11940 20347 11942
rect 20371 11940 20427 11942
rect 20131 10906 20187 10908
rect 20211 10906 20267 10908
rect 20291 10906 20347 10908
rect 20371 10906 20427 10908
rect 20131 10854 20177 10906
rect 20177 10854 20187 10906
rect 20211 10854 20241 10906
rect 20241 10854 20253 10906
rect 20253 10854 20267 10906
rect 20291 10854 20305 10906
rect 20305 10854 20317 10906
rect 20317 10854 20347 10906
rect 20371 10854 20381 10906
rect 20381 10854 20427 10906
rect 20131 10852 20187 10854
rect 20211 10852 20267 10854
rect 20291 10852 20347 10854
rect 20371 10852 20427 10854
rect 20131 9818 20187 9820
rect 20211 9818 20267 9820
rect 20291 9818 20347 9820
rect 20371 9818 20427 9820
rect 20131 9766 20177 9818
rect 20177 9766 20187 9818
rect 20211 9766 20241 9818
rect 20241 9766 20253 9818
rect 20253 9766 20267 9818
rect 20291 9766 20305 9818
rect 20305 9766 20317 9818
rect 20317 9766 20347 9818
rect 20371 9766 20381 9818
rect 20381 9766 20427 9818
rect 20131 9764 20187 9766
rect 20211 9764 20267 9766
rect 20291 9764 20347 9766
rect 20371 9764 20427 9766
rect 22190 11636 22192 11656
rect 22192 11636 22244 11656
rect 22244 11636 22246 11656
rect 22190 11600 22246 11636
rect 20131 8730 20187 8732
rect 20211 8730 20267 8732
rect 20291 8730 20347 8732
rect 20371 8730 20427 8732
rect 20131 8678 20177 8730
rect 20177 8678 20187 8730
rect 20211 8678 20241 8730
rect 20241 8678 20253 8730
rect 20253 8678 20267 8730
rect 20291 8678 20305 8730
rect 20305 8678 20317 8730
rect 20317 8678 20347 8730
rect 20371 8678 20381 8730
rect 20381 8678 20427 8730
rect 20131 8676 20187 8678
rect 20211 8676 20267 8678
rect 20291 8676 20347 8678
rect 20371 8676 20427 8678
rect 19471 8186 19527 8188
rect 19551 8186 19607 8188
rect 19631 8186 19687 8188
rect 19711 8186 19767 8188
rect 19471 8134 19517 8186
rect 19517 8134 19527 8186
rect 19551 8134 19581 8186
rect 19581 8134 19593 8186
rect 19593 8134 19607 8186
rect 19631 8134 19645 8186
rect 19645 8134 19657 8186
rect 19657 8134 19687 8186
rect 19711 8134 19721 8186
rect 19721 8134 19767 8186
rect 19471 8132 19527 8134
rect 19551 8132 19607 8134
rect 19631 8132 19687 8134
rect 19711 8132 19767 8134
rect 14181 3834 14237 3836
rect 14261 3834 14317 3836
rect 14341 3834 14397 3836
rect 14421 3834 14477 3836
rect 14181 3782 14227 3834
rect 14227 3782 14237 3834
rect 14261 3782 14291 3834
rect 14291 3782 14303 3834
rect 14303 3782 14317 3834
rect 14341 3782 14355 3834
rect 14355 3782 14367 3834
rect 14367 3782 14397 3834
rect 14421 3782 14431 3834
rect 14431 3782 14477 3834
rect 14181 3780 14237 3782
rect 14261 3780 14317 3782
rect 14341 3780 14397 3782
rect 14421 3780 14477 3782
rect 3601 2746 3657 2748
rect 3681 2746 3737 2748
rect 3761 2746 3817 2748
rect 3841 2746 3897 2748
rect 3601 2694 3647 2746
rect 3647 2694 3657 2746
rect 3681 2694 3711 2746
rect 3711 2694 3723 2746
rect 3723 2694 3737 2746
rect 3761 2694 3775 2746
rect 3775 2694 3787 2746
rect 3787 2694 3817 2746
rect 3841 2694 3851 2746
rect 3851 2694 3897 2746
rect 3601 2692 3657 2694
rect 3681 2692 3737 2694
rect 3761 2692 3817 2694
rect 3841 2692 3897 2694
rect 8891 2746 8947 2748
rect 8971 2746 9027 2748
rect 9051 2746 9107 2748
rect 9131 2746 9187 2748
rect 8891 2694 8937 2746
rect 8937 2694 8947 2746
rect 8971 2694 9001 2746
rect 9001 2694 9013 2746
rect 9013 2694 9027 2746
rect 9051 2694 9065 2746
rect 9065 2694 9077 2746
rect 9077 2694 9107 2746
rect 9131 2694 9141 2746
rect 9141 2694 9187 2746
rect 8891 2692 8947 2694
rect 8971 2692 9027 2694
rect 9051 2692 9107 2694
rect 9131 2692 9187 2694
rect 14841 3290 14897 3292
rect 14921 3290 14977 3292
rect 15001 3290 15057 3292
rect 15081 3290 15137 3292
rect 14841 3238 14887 3290
rect 14887 3238 14897 3290
rect 14921 3238 14951 3290
rect 14951 3238 14963 3290
rect 14963 3238 14977 3290
rect 15001 3238 15015 3290
rect 15015 3238 15027 3290
rect 15027 3238 15057 3290
rect 15081 3238 15091 3290
rect 15091 3238 15137 3290
rect 14841 3236 14897 3238
rect 14921 3236 14977 3238
rect 15001 3236 15057 3238
rect 15081 3236 15137 3238
rect 14181 2746 14237 2748
rect 14261 2746 14317 2748
rect 14341 2746 14397 2748
rect 14421 2746 14477 2748
rect 14181 2694 14227 2746
rect 14227 2694 14237 2746
rect 14261 2694 14291 2746
rect 14291 2694 14303 2746
rect 14303 2694 14317 2746
rect 14341 2694 14355 2746
rect 14355 2694 14367 2746
rect 14367 2694 14397 2746
rect 14421 2694 14431 2746
rect 14431 2694 14477 2746
rect 14181 2692 14237 2694
rect 14261 2692 14317 2694
rect 14341 2692 14397 2694
rect 14421 2692 14477 2694
rect 20131 7642 20187 7644
rect 20211 7642 20267 7644
rect 20291 7642 20347 7644
rect 20371 7642 20427 7644
rect 20131 7590 20177 7642
rect 20177 7590 20187 7642
rect 20211 7590 20241 7642
rect 20241 7590 20253 7642
rect 20253 7590 20267 7642
rect 20291 7590 20305 7642
rect 20305 7590 20317 7642
rect 20317 7590 20347 7642
rect 20371 7590 20381 7642
rect 20381 7590 20427 7642
rect 20131 7588 20187 7590
rect 20211 7588 20267 7590
rect 20291 7588 20347 7590
rect 20371 7588 20427 7590
rect 19471 7098 19527 7100
rect 19551 7098 19607 7100
rect 19631 7098 19687 7100
rect 19711 7098 19767 7100
rect 19471 7046 19517 7098
rect 19517 7046 19527 7098
rect 19551 7046 19581 7098
rect 19581 7046 19593 7098
rect 19593 7046 19607 7098
rect 19631 7046 19645 7098
rect 19645 7046 19657 7098
rect 19657 7046 19687 7098
rect 19711 7046 19721 7098
rect 19721 7046 19767 7098
rect 19471 7044 19527 7046
rect 19551 7044 19607 7046
rect 19631 7044 19687 7046
rect 19711 7044 19767 7046
rect 20131 6554 20187 6556
rect 20211 6554 20267 6556
rect 20291 6554 20347 6556
rect 20371 6554 20427 6556
rect 20131 6502 20177 6554
rect 20177 6502 20187 6554
rect 20211 6502 20241 6554
rect 20241 6502 20253 6554
rect 20253 6502 20267 6554
rect 20291 6502 20305 6554
rect 20305 6502 20317 6554
rect 20317 6502 20347 6554
rect 20371 6502 20381 6554
rect 20381 6502 20427 6554
rect 20131 6500 20187 6502
rect 20211 6500 20267 6502
rect 20291 6500 20347 6502
rect 20371 6500 20427 6502
rect 19471 6010 19527 6012
rect 19551 6010 19607 6012
rect 19631 6010 19687 6012
rect 19711 6010 19767 6012
rect 19471 5958 19517 6010
rect 19517 5958 19527 6010
rect 19551 5958 19581 6010
rect 19581 5958 19593 6010
rect 19593 5958 19607 6010
rect 19631 5958 19645 6010
rect 19645 5958 19657 6010
rect 19657 5958 19687 6010
rect 19711 5958 19721 6010
rect 19721 5958 19767 6010
rect 19471 5956 19527 5958
rect 19551 5956 19607 5958
rect 19631 5956 19687 5958
rect 19711 5956 19767 5958
rect 20131 5466 20187 5468
rect 20211 5466 20267 5468
rect 20291 5466 20347 5468
rect 20371 5466 20427 5468
rect 20131 5414 20177 5466
rect 20177 5414 20187 5466
rect 20211 5414 20241 5466
rect 20241 5414 20253 5466
rect 20253 5414 20267 5466
rect 20291 5414 20305 5466
rect 20305 5414 20317 5466
rect 20317 5414 20347 5466
rect 20371 5414 20381 5466
rect 20381 5414 20427 5466
rect 20131 5412 20187 5414
rect 20211 5412 20267 5414
rect 20291 5412 20347 5414
rect 20371 5412 20427 5414
rect 19471 4922 19527 4924
rect 19551 4922 19607 4924
rect 19631 4922 19687 4924
rect 19711 4922 19767 4924
rect 19471 4870 19517 4922
rect 19517 4870 19527 4922
rect 19551 4870 19581 4922
rect 19581 4870 19593 4922
rect 19593 4870 19607 4922
rect 19631 4870 19645 4922
rect 19645 4870 19657 4922
rect 19657 4870 19687 4922
rect 19711 4870 19721 4922
rect 19721 4870 19767 4922
rect 19471 4868 19527 4870
rect 19551 4868 19607 4870
rect 19631 4868 19687 4870
rect 19711 4868 19767 4870
rect 20131 4378 20187 4380
rect 20211 4378 20267 4380
rect 20291 4378 20347 4380
rect 20371 4378 20427 4380
rect 20131 4326 20177 4378
rect 20177 4326 20187 4378
rect 20211 4326 20241 4378
rect 20241 4326 20253 4378
rect 20253 4326 20267 4378
rect 20291 4326 20305 4378
rect 20305 4326 20317 4378
rect 20317 4326 20347 4378
rect 20371 4326 20381 4378
rect 20381 4326 20427 4378
rect 20131 4324 20187 4326
rect 20211 4324 20267 4326
rect 20291 4324 20347 4326
rect 20371 4324 20427 4326
rect 19471 3834 19527 3836
rect 19551 3834 19607 3836
rect 19631 3834 19687 3836
rect 19711 3834 19767 3836
rect 19471 3782 19517 3834
rect 19517 3782 19527 3834
rect 19551 3782 19581 3834
rect 19581 3782 19593 3834
rect 19593 3782 19607 3834
rect 19631 3782 19645 3834
rect 19645 3782 19657 3834
rect 19657 3782 19687 3834
rect 19711 3782 19721 3834
rect 19721 3782 19767 3834
rect 19471 3780 19527 3782
rect 19551 3780 19607 3782
rect 19631 3780 19687 3782
rect 19711 3780 19767 3782
rect 20131 3290 20187 3292
rect 20211 3290 20267 3292
rect 20291 3290 20347 3292
rect 20371 3290 20427 3292
rect 20131 3238 20177 3290
rect 20177 3238 20187 3290
rect 20211 3238 20241 3290
rect 20241 3238 20253 3290
rect 20253 3238 20267 3290
rect 20291 3238 20305 3290
rect 20305 3238 20317 3290
rect 20317 3238 20347 3290
rect 20371 3238 20381 3290
rect 20381 3238 20427 3290
rect 20131 3236 20187 3238
rect 20211 3236 20267 3238
rect 20291 3236 20347 3238
rect 20371 3236 20427 3238
rect 19471 2746 19527 2748
rect 19551 2746 19607 2748
rect 19631 2746 19687 2748
rect 19711 2746 19767 2748
rect 19471 2694 19517 2746
rect 19517 2694 19527 2746
rect 19551 2694 19581 2746
rect 19581 2694 19593 2746
rect 19593 2694 19607 2746
rect 19631 2694 19645 2746
rect 19645 2694 19657 2746
rect 19657 2694 19687 2746
rect 19711 2694 19721 2746
rect 19721 2694 19767 2746
rect 19471 2692 19527 2694
rect 19551 2692 19607 2694
rect 19631 2692 19687 2694
rect 19711 2692 19767 2694
rect 4261 2202 4317 2204
rect 4341 2202 4397 2204
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4261 2150 4307 2202
rect 4307 2150 4317 2202
rect 4341 2150 4371 2202
rect 4371 2150 4383 2202
rect 4383 2150 4397 2202
rect 4421 2150 4435 2202
rect 4435 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4261 2148 4317 2150
rect 4341 2148 4397 2150
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 9551 2202 9607 2204
rect 9631 2202 9687 2204
rect 9711 2202 9767 2204
rect 9791 2202 9847 2204
rect 9551 2150 9597 2202
rect 9597 2150 9607 2202
rect 9631 2150 9661 2202
rect 9661 2150 9673 2202
rect 9673 2150 9687 2202
rect 9711 2150 9725 2202
rect 9725 2150 9737 2202
rect 9737 2150 9767 2202
rect 9791 2150 9801 2202
rect 9801 2150 9847 2202
rect 9551 2148 9607 2150
rect 9631 2148 9687 2150
rect 9711 2148 9767 2150
rect 9791 2148 9847 2150
rect 14841 2202 14897 2204
rect 14921 2202 14977 2204
rect 15001 2202 15057 2204
rect 15081 2202 15137 2204
rect 14841 2150 14887 2202
rect 14887 2150 14897 2202
rect 14921 2150 14951 2202
rect 14951 2150 14963 2202
rect 14963 2150 14977 2202
rect 15001 2150 15015 2202
rect 15015 2150 15027 2202
rect 15027 2150 15057 2202
rect 15081 2150 15091 2202
rect 15091 2150 15137 2202
rect 14841 2148 14897 2150
rect 14921 2148 14977 2150
rect 15001 2148 15057 2150
rect 15081 2148 15137 2150
rect 20131 2202 20187 2204
rect 20211 2202 20267 2204
rect 20291 2202 20347 2204
rect 20371 2202 20427 2204
rect 20131 2150 20177 2202
rect 20177 2150 20187 2202
rect 20211 2150 20241 2202
rect 20241 2150 20253 2202
rect 20253 2150 20267 2202
rect 20291 2150 20305 2202
rect 20305 2150 20317 2202
rect 20317 2150 20347 2202
rect 20371 2150 20381 2202
rect 20381 2150 20427 2202
rect 20131 2148 20187 2150
rect 20211 2148 20267 2150
rect 20291 2148 20347 2150
rect 20371 2148 20427 2150
rect 22190 2080 22246 2136
<< metal3 >>
rect 4251 22880 4567 22881
rect 4251 22816 4257 22880
rect 4321 22816 4337 22880
rect 4401 22816 4417 22880
rect 4481 22816 4497 22880
rect 4561 22816 4567 22880
rect 4251 22815 4567 22816
rect 9541 22880 9857 22881
rect 9541 22816 9547 22880
rect 9611 22816 9627 22880
rect 9691 22816 9707 22880
rect 9771 22816 9787 22880
rect 9851 22816 9857 22880
rect 9541 22815 9857 22816
rect 14831 22880 15147 22881
rect 14831 22816 14837 22880
rect 14901 22816 14917 22880
rect 14981 22816 14997 22880
rect 15061 22816 15077 22880
rect 15141 22816 15147 22880
rect 14831 22815 15147 22816
rect 20121 22880 20437 22881
rect 20121 22816 20127 22880
rect 20191 22816 20207 22880
rect 20271 22816 20287 22880
rect 20351 22816 20367 22880
rect 20431 22816 20437 22880
rect 20121 22815 20437 22816
rect 3591 22336 3907 22337
rect 3591 22272 3597 22336
rect 3661 22272 3677 22336
rect 3741 22272 3757 22336
rect 3821 22272 3837 22336
rect 3901 22272 3907 22336
rect 3591 22271 3907 22272
rect 8881 22336 9197 22337
rect 8881 22272 8887 22336
rect 8951 22272 8967 22336
rect 9031 22272 9047 22336
rect 9111 22272 9127 22336
rect 9191 22272 9197 22336
rect 8881 22271 9197 22272
rect 14171 22336 14487 22337
rect 14171 22272 14177 22336
rect 14241 22272 14257 22336
rect 14321 22272 14337 22336
rect 14401 22272 14417 22336
rect 14481 22272 14487 22336
rect 14171 22271 14487 22272
rect 19461 22336 19777 22337
rect 19461 22272 19467 22336
rect 19531 22272 19547 22336
rect 19611 22272 19627 22336
rect 19691 22272 19707 22336
rect 19771 22272 19777 22336
rect 19461 22271 19777 22272
rect 4251 21792 4567 21793
rect 4251 21728 4257 21792
rect 4321 21728 4337 21792
rect 4401 21728 4417 21792
rect 4481 21728 4497 21792
rect 4561 21728 4567 21792
rect 4251 21727 4567 21728
rect 9541 21792 9857 21793
rect 9541 21728 9547 21792
rect 9611 21728 9627 21792
rect 9691 21728 9707 21792
rect 9771 21728 9787 21792
rect 9851 21728 9857 21792
rect 9541 21727 9857 21728
rect 14831 21792 15147 21793
rect 14831 21728 14837 21792
rect 14901 21728 14917 21792
rect 14981 21728 14997 21792
rect 15061 21728 15077 21792
rect 15141 21728 15147 21792
rect 14831 21727 15147 21728
rect 20121 21792 20437 21793
rect 20121 21728 20127 21792
rect 20191 21728 20207 21792
rect 20271 21728 20287 21792
rect 20351 21728 20367 21792
rect 20431 21728 20437 21792
rect 20121 21727 20437 21728
rect 6729 21450 6795 21453
rect 7649 21450 7715 21453
rect 6729 21448 7715 21450
rect 6729 21392 6734 21448
rect 6790 21392 7654 21448
rect 7710 21392 7715 21448
rect 6729 21390 7715 21392
rect 6729 21387 6795 21390
rect 7649 21387 7715 21390
rect 16297 21314 16363 21317
rect 16941 21314 17007 21317
rect 16297 21312 17007 21314
rect 16297 21256 16302 21312
rect 16358 21256 16946 21312
rect 17002 21256 17007 21312
rect 16297 21254 17007 21256
rect 16297 21251 16363 21254
rect 16941 21251 17007 21254
rect 3591 21248 3907 21249
rect 3591 21184 3597 21248
rect 3661 21184 3677 21248
rect 3741 21184 3757 21248
rect 3821 21184 3837 21248
rect 3901 21184 3907 21248
rect 3591 21183 3907 21184
rect 8881 21248 9197 21249
rect 8881 21184 8887 21248
rect 8951 21184 8967 21248
rect 9031 21184 9047 21248
rect 9111 21184 9127 21248
rect 9191 21184 9197 21248
rect 8881 21183 9197 21184
rect 14171 21248 14487 21249
rect 14171 21184 14177 21248
rect 14241 21184 14257 21248
rect 14321 21184 14337 21248
rect 14401 21184 14417 21248
rect 14481 21184 14487 21248
rect 14171 21183 14487 21184
rect 19461 21248 19777 21249
rect 19461 21184 19467 21248
rect 19531 21184 19547 21248
rect 19611 21184 19627 21248
rect 19691 21184 19707 21248
rect 19771 21184 19777 21248
rect 19461 21183 19777 21184
rect 22185 21178 22251 21181
rect 22608 21178 23408 21208
rect 22185 21176 23408 21178
rect 22185 21120 22190 21176
rect 22246 21120 23408 21176
rect 22185 21118 23408 21120
rect 22185 21115 22251 21118
rect 22608 21088 23408 21118
rect 4251 20704 4567 20705
rect 4251 20640 4257 20704
rect 4321 20640 4337 20704
rect 4401 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4567 20704
rect 4251 20639 4567 20640
rect 9541 20704 9857 20705
rect 9541 20640 9547 20704
rect 9611 20640 9627 20704
rect 9691 20640 9707 20704
rect 9771 20640 9787 20704
rect 9851 20640 9857 20704
rect 9541 20639 9857 20640
rect 14831 20704 15147 20705
rect 14831 20640 14837 20704
rect 14901 20640 14917 20704
rect 14981 20640 14997 20704
rect 15061 20640 15077 20704
rect 15141 20640 15147 20704
rect 14831 20639 15147 20640
rect 20121 20704 20437 20705
rect 20121 20640 20127 20704
rect 20191 20640 20207 20704
rect 20271 20640 20287 20704
rect 20351 20640 20367 20704
rect 20431 20640 20437 20704
rect 20121 20639 20437 20640
rect 3591 20160 3907 20161
rect 3591 20096 3597 20160
rect 3661 20096 3677 20160
rect 3741 20096 3757 20160
rect 3821 20096 3837 20160
rect 3901 20096 3907 20160
rect 3591 20095 3907 20096
rect 8881 20160 9197 20161
rect 8881 20096 8887 20160
rect 8951 20096 8967 20160
rect 9031 20096 9047 20160
rect 9111 20096 9127 20160
rect 9191 20096 9197 20160
rect 8881 20095 9197 20096
rect 14171 20160 14487 20161
rect 14171 20096 14177 20160
rect 14241 20096 14257 20160
rect 14321 20096 14337 20160
rect 14401 20096 14417 20160
rect 14481 20096 14487 20160
rect 14171 20095 14487 20096
rect 19461 20160 19777 20161
rect 19461 20096 19467 20160
rect 19531 20096 19547 20160
rect 19611 20096 19627 20160
rect 19691 20096 19707 20160
rect 19771 20096 19777 20160
rect 19461 20095 19777 20096
rect 4251 19616 4567 19617
rect 4251 19552 4257 19616
rect 4321 19552 4337 19616
rect 4401 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4567 19616
rect 4251 19551 4567 19552
rect 9541 19616 9857 19617
rect 9541 19552 9547 19616
rect 9611 19552 9627 19616
rect 9691 19552 9707 19616
rect 9771 19552 9787 19616
rect 9851 19552 9857 19616
rect 9541 19551 9857 19552
rect 14831 19616 15147 19617
rect 14831 19552 14837 19616
rect 14901 19552 14917 19616
rect 14981 19552 14997 19616
rect 15061 19552 15077 19616
rect 15141 19552 15147 19616
rect 14831 19551 15147 19552
rect 20121 19616 20437 19617
rect 20121 19552 20127 19616
rect 20191 19552 20207 19616
rect 20271 19552 20287 19616
rect 20351 19552 20367 19616
rect 20431 19552 20437 19616
rect 20121 19551 20437 19552
rect 11329 19410 11395 19413
rect 12157 19410 12223 19413
rect 16573 19410 16639 19413
rect 11329 19408 16639 19410
rect 11329 19352 11334 19408
rect 11390 19352 12162 19408
rect 12218 19352 16578 19408
rect 16634 19352 16639 19408
rect 11329 19350 16639 19352
rect 11329 19347 11395 19350
rect 12157 19347 12223 19350
rect 16573 19347 16639 19350
rect 3591 19072 3907 19073
rect 3591 19008 3597 19072
rect 3661 19008 3677 19072
rect 3741 19008 3757 19072
rect 3821 19008 3837 19072
rect 3901 19008 3907 19072
rect 3591 19007 3907 19008
rect 8881 19072 9197 19073
rect 8881 19008 8887 19072
rect 8951 19008 8967 19072
rect 9031 19008 9047 19072
rect 9111 19008 9127 19072
rect 9191 19008 9197 19072
rect 8881 19007 9197 19008
rect 14171 19072 14487 19073
rect 14171 19008 14177 19072
rect 14241 19008 14257 19072
rect 14321 19008 14337 19072
rect 14401 19008 14417 19072
rect 14481 19008 14487 19072
rect 14171 19007 14487 19008
rect 19461 19072 19777 19073
rect 19461 19008 19467 19072
rect 19531 19008 19547 19072
rect 19611 19008 19627 19072
rect 19691 19008 19707 19072
rect 19771 19008 19777 19072
rect 19461 19007 19777 19008
rect 4251 18528 4567 18529
rect 0 18458 800 18488
rect 4251 18464 4257 18528
rect 4321 18464 4337 18528
rect 4401 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4567 18528
rect 4251 18463 4567 18464
rect 9541 18528 9857 18529
rect 9541 18464 9547 18528
rect 9611 18464 9627 18528
rect 9691 18464 9707 18528
rect 9771 18464 9787 18528
rect 9851 18464 9857 18528
rect 9541 18463 9857 18464
rect 14831 18528 15147 18529
rect 14831 18464 14837 18528
rect 14901 18464 14917 18528
rect 14981 18464 14997 18528
rect 15061 18464 15077 18528
rect 15141 18464 15147 18528
rect 14831 18463 15147 18464
rect 20121 18528 20437 18529
rect 20121 18464 20127 18528
rect 20191 18464 20207 18528
rect 20271 18464 20287 18528
rect 20351 18464 20367 18528
rect 20431 18464 20437 18528
rect 20121 18463 20437 18464
rect 5073 18458 5139 18461
rect 0 18398 4170 18458
rect 0 18368 800 18398
rect 4110 18322 4170 18398
rect 4662 18456 5139 18458
rect 4662 18400 5078 18456
rect 5134 18400 5139 18456
rect 4662 18398 5139 18400
rect 4662 18322 4722 18398
rect 5073 18395 5139 18398
rect 4110 18262 4722 18322
rect 13997 18186 14063 18189
rect 15561 18186 15627 18189
rect 13997 18184 15627 18186
rect 13997 18128 14002 18184
rect 14058 18128 15566 18184
rect 15622 18128 15627 18184
rect 13997 18126 15627 18128
rect 13997 18123 14063 18126
rect 15561 18123 15627 18126
rect 3591 17984 3907 17985
rect 3591 17920 3597 17984
rect 3661 17920 3677 17984
rect 3741 17920 3757 17984
rect 3821 17920 3837 17984
rect 3901 17920 3907 17984
rect 3591 17919 3907 17920
rect 8881 17984 9197 17985
rect 8881 17920 8887 17984
rect 8951 17920 8967 17984
rect 9031 17920 9047 17984
rect 9111 17920 9127 17984
rect 9191 17920 9197 17984
rect 8881 17919 9197 17920
rect 14171 17984 14487 17985
rect 14171 17920 14177 17984
rect 14241 17920 14257 17984
rect 14321 17920 14337 17984
rect 14401 17920 14417 17984
rect 14481 17920 14487 17984
rect 14171 17919 14487 17920
rect 19461 17984 19777 17985
rect 19461 17920 19467 17984
rect 19531 17920 19547 17984
rect 19611 17920 19627 17984
rect 19691 17920 19707 17984
rect 19771 17920 19777 17984
rect 19461 17919 19777 17920
rect 4251 17440 4567 17441
rect 4251 17376 4257 17440
rect 4321 17376 4337 17440
rect 4401 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4567 17440
rect 4251 17375 4567 17376
rect 9541 17440 9857 17441
rect 9541 17376 9547 17440
rect 9611 17376 9627 17440
rect 9691 17376 9707 17440
rect 9771 17376 9787 17440
rect 9851 17376 9857 17440
rect 9541 17375 9857 17376
rect 14831 17440 15147 17441
rect 14831 17376 14837 17440
rect 14901 17376 14917 17440
rect 14981 17376 14997 17440
rect 15061 17376 15077 17440
rect 15141 17376 15147 17440
rect 14831 17375 15147 17376
rect 20121 17440 20437 17441
rect 20121 17376 20127 17440
rect 20191 17376 20207 17440
rect 20271 17376 20287 17440
rect 20351 17376 20367 17440
rect 20431 17376 20437 17440
rect 20121 17375 20437 17376
rect 9213 17234 9279 17237
rect 9489 17234 9555 17237
rect 9213 17232 9555 17234
rect 9213 17176 9218 17232
rect 9274 17176 9494 17232
rect 9550 17176 9555 17232
rect 9213 17174 9555 17176
rect 9213 17171 9279 17174
rect 9489 17171 9555 17174
rect 3591 16896 3907 16897
rect 3591 16832 3597 16896
rect 3661 16832 3677 16896
rect 3741 16832 3757 16896
rect 3821 16832 3837 16896
rect 3901 16832 3907 16896
rect 3591 16831 3907 16832
rect 8881 16896 9197 16897
rect 8881 16832 8887 16896
rect 8951 16832 8967 16896
rect 9031 16832 9047 16896
rect 9111 16832 9127 16896
rect 9191 16832 9197 16896
rect 8881 16831 9197 16832
rect 14171 16896 14487 16897
rect 14171 16832 14177 16896
rect 14241 16832 14257 16896
rect 14321 16832 14337 16896
rect 14401 16832 14417 16896
rect 14481 16832 14487 16896
rect 14171 16831 14487 16832
rect 19461 16896 19777 16897
rect 19461 16832 19467 16896
rect 19531 16832 19547 16896
rect 19611 16832 19627 16896
rect 19691 16832 19707 16896
rect 19771 16832 19777 16896
rect 19461 16831 19777 16832
rect 20069 16554 20135 16557
rect 19934 16552 20135 16554
rect 19934 16496 20074 16552
rect 20130 16496 20135 16552
rect 19934 16494 20135 16496
rect 4251 16352 4567 16353
rect 4251 16288 4257 16352
rect 4321 16288 4337 16352
rect 4401 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4567 16352
rect 4251 16287 4567 16288
rect 9541 16352 9857 16353
rect 9541 16288 9547 16352
rect 9611 16288 9627 16352
rect 9691 16288 9707 16352
rect 9771 16288 9787 16352
rect 9851 16288 9857 16352
rect 9541 16287 9857 16288
rect 14831 16352 15147 16353
rect 14831 16288 14837 16352
rect 14901 16288 14917 16352
rect 14981 16288 14997 16352
rect 15061 16288 15077 16352
rect 15141 16288 15147 16352
rect 14831 16287 15147 16288
rect 19934 16149 19994 16494
rect 20069 16491 20135 16494
rect 20121 16352 20437 16353
rect 20121 16288 20127 16352
rect 20191 16288 20207 16352
rect 20271 16288 20287 16352
rect 20351 16288 20367 16352
rect 20431 16288 20437 16352
rect 20121 16287 20437 16288
rect 19934 16144 20043 16149
rect 19934 16088 19982 16144
rect 20038 16088 20043 16144
rect 19934 16086 20043 16088
rect 19977 16083 20043 16086
rect 19609 16010 19675 16013
rect 19609 16008 19994 16010
rect 19609 15952 19614 16008
rect 19670 15952 19994 16008
rect 19609 15950 19994 15952
rect 19609 15947 19675 15950
rect 3591 15808 3907 15809
rect 3591 15744 3597 15808
rect 3661 15744 3677 15808
rect 3741 15744 3757 15808
rect 3821 15744 3837 15808
rect 3901 15744 3907 15808
rect 3591 15743 3907 15744
rect 8881 15808 9197 15809
rect 8881 15744 8887 15808
rect 8951 15744 8967 15808
rect 9031 15744 9047 15808
rect 9111 15744 9127 15808
rect 9191 15744 9197 15808
rect 8881 15743 9197 15744
rect 14171 15808 14487 15809
rect 14171 15744 14177 15808
rect 14241 15744 14257 15808
rect 14321 15744 14337 15808
rect 14401 15744 14417 15808
rect 14481 15744 14487 15808
rect 14171 15743 14487 15744
rect 19461 15808 19777 15809
rect 19461 15744 19467 15808
rect 19531 15744 19547 15808
rect 19611 15744 19627 15808
rect 19691 15744 19707 15808
rect 19771 15744 19777 15808
rect 19461 15743 19777 15744
rect 11881 15602 11947 15605
rect 15285 15602 15351 15605
rect 11881 15600 15351 15602
rect 11881 15544 11886 15600
rect 11942 15544 15290 15600
rect 15346 15544 15351 15600
rect 11881 15542 15351 15544
rect 11881 15539 11947 15542
rect 15285 15539 15351 15542
rect 19333 15602 19399 15605
rect 19934 15602 19994 15950
rect 19333 15600 19994 15602
rect 19333 15544 19338 15600
rect 19394 15544 19994 15600
rect 19333 15542 19994 15544
rect 19333 15539 19399 15542
rect 4251 15264 4567 15265
rect 4251 15200 4257 15264
rect 4321 15200 4337 15264
rect 4401 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4567 15264
rect 4251 15199 4567 15200
rect 9541 15264 9857 15265
rect 9541 15200 9547 15264
rect 9611 15200 9627 15264
rect 9691 15200 9707 15264
rect 9771 15200 9787 15264
rect 9851 15200 9857 15264
rect 9541 15199 9857 15200
rect 14831 15264 15147 15265
rect 14831 15200 14837 15264
rect 14901 15200 14917 15264
rect 14981 15200 14997 15264
rect 15061 15200 15077 15264
rect 15141 15200 15147 15264
rect 14831 15199 15147 15200
rect 20121 15264 20437 15265
rect 20121 15200 20127 15264
rect 20191 15200 20207 15264
rect 20271 15200 20287 15264
rect 20351 15200 20367 15264
rect 20431 15200 20437 15264
rect 20121 15199 20437 15200
rect 3591 14720 3907 14721
rect 3591 14656 3597 14720
rect 3661 14656 3677 14720
rect 3741 14656 3757 14720
rect 3821 14656 3837 14720
rect 3901 14656 3907 14720
rect 3591 14655 3907 14656
rect 8881 14720 9197 14721
rect 8881 14656 8887 14720
rect 8951 14656 8967 14720
rect 9031 14656 9047 14720
rect 9111 14656 9127 14720
rect 9191 14656 9197 14720
rect 8881 14655 9197 14656
rect 14171 14720 14487 14721
rect 14171 14656 14177 14720
rect 14241 14656 14257 14720
rect 14321 14656 14337 14720
rect 14401 14656 14417 14720
rect 14481 14656 14487 14720
rect 14171 14655 14487 14656
rect 19461 14720 19777 14721
rect 19461 14656 19467 14720
rect 19531 14656 19547 14720
rect 19611 14656 19627 14720
rect 19691 14656 19707 14720
rect 19771 14656 19777 14720
rect 19461 14655 19777 14656
rect 4251 14176 4567 14177
rect 4251 14112 4257 14176
rect 4321 14112 4337 14176
rect 4401 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4567 14176
rect 4251 14111 4567 14112
rect 9541 14176 9857 14177
rect 9541 14112 9547 14176
rect 9611 14112 9627 14176
rect 9691 14112 9707 14176
rect 9771 14112 9787 14176
rect 9851 14112 9857 14176
rect 9541 14111 9857 14112
rect 14831 14176 15147 14177
rect 14831 14112 14837 14176
rect 14901 14112 14917 14176
rect 14981 14112 14997 14176
rect 15061 14112 15077 14176
rect 15141 14112 15147 14176
rect 14831 14111 15147 14112
rect 20121 14176 20437 14177
rect 20121 14112 20127 14176
rect 20191 14112 20207 14176
rect 20271 14112 20287 14176
rect 20351 14112 20367 14176
rect 20431 14112 20437 14176
rect 20121 14111 20437 14112
rect 3591 13632 3907 13633
rect 3591 13568 3597 13632
rect 3661 13568 3677 13632
rect 3741 13568 3757 13632
rect 3821 13568 3837 13632
rect 3901 13568 3907 13632
rect 3591 13567 3907 13568
rect 8881 13632 9197 13633
rect 8881 13568 8887 13632
rect 8951 13568 8967 13632
rect 9031 13568 9047 13632
rect 9111 13568 9127 13632
rect 9191 13568 9197 13632
rect 8881 13567 9197 13568
rect 14171 13632 14487 13633
rect 14171 13568 14177 13632
rect 14241 13568 14257 13632
rect 14321 13568 14337 13632
rect 14401 13568 14417 13632
rect 14481 13568 14487 13632
rect 14171 13567 14487 13568
rect 19461 13632 19777 13633
rect 19461 13568 19467 13632
rect 19531 13568 19547 13632
rect 19611 13568 19627 13632
rect 19691 13568 19707 13632
rect 19771 13568 19777 13632
rect 19461 13567 19777 13568
rect 4251 13088 4567 13089
rect 4251 13024 4257 13088
rect 4321 13024 4337 13088
rect 4401 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4567 13088
rect 4251 13023 4567 13024
rect 9541 13088 9857 13089
rect 9541 13024 9547 13088
rect 9611 13024 9627 13088
rect 9691 13024 9707 13088
rect 9771 13024 9787 13088
rect 9851 13024 9857 13088
rect 9541 13023 9857 13024
rect 14831 13088 15147 13089
rect 14831 13024 14837 13088
rect 14901 13024 14917 13088
rect 14981 13024 14997 13088
rect 15061 13024 15077 13088
rect 15141 13024 15147 13088
rect 14831 13023 15147 13024
rect 20121 13088 20437 13089
rect 20121 13024 20127 13088
rect 20191 13024 20207 13088
rect 20271 13024 20287 13088
rect 20351 13024 20367 13088
rect 20431 13024 20437 13088
rect 20121 13023 20437 13024
rect 3591 12544 3907 12545
rect 3591 12480 3597 12544
rect 3661 12480 3677 12544
rect 3741 12480 3757 12544
rect 3821 12480 3837 12544
rect 3901 12480 3907 12544
rect 3591 12479 3907 12480
rect 8881 12544 9197 12545
rect 8881 12480 8887 12544
rect 8951 12480 8967 12544
rect 9031 12480 9047 12544
rect 9111 12480 9127 12544
rect 9191 12480 9197 12544
rect 8881 12479 9197 12480
rect 14171 12544 14487 12545
rect 14171 12480 14177 12544
rect 14241 12480 14257 12544
rect 14321 12480 14337 12544
rect 14401 12480 14417 12544
rect 14481 12480 14487 12544
rect 14171 12479 14487 12480
rect 19461 12544 19777 12545
rect 19461 12480 19467 12544
rect 19531 12480 19547 12544
rect 19611 12480 19627 12544
rect 19691 12480 19707 12544
rect 19771 12480 19777 12544
rect 19461 12479 19777 12480
rect 4251 12000 4567 12001
rect 4251 11936 4257 12000
rect 4321 11936 4337 12000
rect 4401 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4567 12000
rect 4251 11935 4567 11936
rect 9541 12000 9857 12001
rect 9541 11936 9547 12000
rect 9611 11936 9627 12000
rect 9691 11936 9707 12000
rect 9771 11936 9787 12000
rect 9851 11936 9857 12000
rect 9541 11935 9857 11936
rect 14831 12000 15147 12001
rect 14831 11936 14837 12000
rect 14901 11936 14917 12000
rect 14981 11936 14997 12000
rect 15061 11936 15077 12000
rect 15141 11936 15147 12000
rect 14831 11935 15147 11936
rect 20121 12000 20437 12001
rect 20121 11936 20127 12000
rect 20191 11936 20207 12000
rect 20271 11936 20287 12000
rect 20351 11936 20367 12000
rect 20431 11936 20437 12000
rect 20121 11935 20437 11936
rect 22185 11658 22251 11661
rect 22608 11658 23408 11688
rect 22185 11656 23408 11658
rect 22185 11600 22190 11656
rect 22246 11600 23408 11656
rect 22185 11598 23408 11600
rect 22185 11595 22251 11598
rect 22608 11568 23408 11598
rect 3591 11456 3907 11457
rect 3591 11392 3597 11456
rect 3661 11392 3677 11456
rect 3741 11392 3757 11456
rect 3821 11392 3837 11456
rect 3901 11392 3907 11456
rect 3591 11391 3907 11392
rect 8881 11456 9197 11457
rect 8881 11392 8887 11456
rect 8951 11392 8967 11456
rect 9031 11392 9047 11456
rect 9111 11392 9127 11456
rect 9191 11392 9197 11456
rect 8881 11391 9197 11392
rect 14171 11456 14487 11457
rect 14171 11392 14177 11456
rect 14241 11392 14257 11456
rect 14321 11392 14337 11456
rect 14401 11392 14417 11456
rect 14481 11392 14487 11456
rect 14171 11391 14487 11392
rect 19461 11456 19777 11457
rect 19461 11392 19467 11456
rect 19531 11392 19547 11456
rect 19611 11392 19627 11456
rect 19691 11392 19707 11456
rect 19771 11392 19777 11456
rect 19461 11391 19777 11392
rect 4251 10912 4567 10913
rect 4251 10848 4257 10912
rect 4321 10848 4337 10912
rect 4401 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4567 10912
rect 4251 10847 4567 10848
rect 9541 10912 9857 10913
rect 9541 10848 9547 10912
rect 9611 10848 9627 10912
rect 9691 10848 9707 10912
rect 9771 10848 9787 10912
rect 9851 10848 9857 10912
rect 9541 10847 9857 10848
rect 14831 10912 15147 10913
rect 14831 10848 14837 10912
rect 14901 10848 14917 10912
rect 14981 10848 14997 10912
rect 15061 10848 15077 10912
rect 15141 10848 15147 10912
rect 14831 10847 15147 10848
rect 20121 10912 20437 10913
rect 20121 10848 20127 10912
rect 20191 10848 20207 10912
rect 20271 10848 20287 10912
rect 20351 10848 20367 10912
rect 20431 10848 20437 10912
rect 20121 10847 20437 10848
rect 3591 10368 3907 10369
rect 3591 10304 3597 10368
rect 3661 10304 3677 10368
rect 3741 10304 3757 10368
rect 3821 10304 3837 10368
rect 3901 10304 3907 10368
rect 3591 10303 3907 10304
rect 8881 10368 9197 10369
rect 8881 10304 8887 10368
rect 8951 10304 8967 10368
rect 9031 10304 9047 10368
rect 9111 10304 9127 10368
rect 9191 10304 9197 10368
rect 8881 10303 9197 10304
rect 14171 10368 14487 10369
rect 14171 10304 14177 10368
rect 14241 10304 14257 10368
rect 14321 10304 14337 10368
rect 14401 10304 14417 10368
rect 14481 10304 14487 10368
rect 14171 10303 14487 10304
rect 19461 10368 19777 10369
rect 19461 10304 19467 10368
rect 19531 10304 19547 10368
rect 19611 10304 19627 10368
rect 19691 10304 19707 10368
rect 19771 10304 19777 10368
rect 19461 10303 19777 10304
rect 4251 9824 4567 9825
rect 4251 9760 4257 9824
rect 4321 9760 4337 9824
rect 4401 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4567 9824
rect 4251 9759 4567 9760
rect 9541 9824 9857 9825
rect 9541 9760 9547 9824
rect 9611 9760 9627 9824
rect 9691 9760 9707 9824
rect 9771 9760 9787 9824
rect 9851 9760 9857 9824
rect 9541 9759 9857 9760
rect 14831 9824 15147 9825
rect 14831 9760 14837 9824
rect 14901 9760 14917 9824
rect 14981 9760 14997 9824
rect 15061 9760 15077 9824
rect 15141 9760 15147 9824
rect 14831 9759 15147 9760
rect 20121 9824 20437 9825
rect 20121 9760 20127 9824
rect 20191 9760 20207 9824
rect 20271 9760 20287 9824
rect 20351 9760 20367 9824
rect 20431 9760 20437 9824
rect 20121 9759 20437 9760
rect 3591 9280 3907 9281
rect 3591 9216 3597 9280
rect 3661 9216 3677 9280
rect 3741 9216 3757 9280
rect 3821 9216 3837 9280
rect 3901 9216 3907 9280
rect 3591 9215 3907 9216
rect 8881 9280 9197 9281
rect 8881 9216 8887 9280
rect 8951 9216 8967 9280
rect 9031 9216 9047 9280
rect 9111 9216 9127 9280
rect 9191 9216 9197 9280
rect 8881 9215 9197 9216
rect 14171 9280 14487 9281
rect 14171 9216 14177 9280
rect 14241 9216 14257 9280
rect 14321 9216 14337 9280
rect 14401 9216 14417 9280
rect 14481 9216 14487 9280
rect 14171 9215 14487 9216
rect 19461 9280 19777 9281
rect 19461 9216 19467 9280
rect 19531 9216 19547 9280
rect 19611 9216 19627 9280
rect 19691 9216 19707 9280
rect 19771 9216 19777 9280
rect 19461 9215 19777 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 4251 8736 4567 8737
rect 4251 8672 4257 8736
rect 4321 8672 4337 8736
rect 4401 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4567 8736
rect 4251 8671 4567 8672
rect 9541 8736 9857 8737
rect 9541 8672 9547 8736
rect 9611 8672 9627 8736
rect 9691 8672 9707 8736
rect 9771 8672 9787 8736
rect 9851 8672 9857 8736
rect 9541 8671 9857 8672
rect 14831 8736 15147 8737
rect 14831 8672 14837 8736
rect 14901 8672 14917 8736
rect 14981 8672 14997 8736
rect 15061 8672 15077 8736
rect 15141 8672 15147 8736
rect 14831 8671 15147 8672
rect 20121 8736 20437 8737
rect 20121 8672 20127 8736
rect 20191 8672 20207 8736
rect 20271 8672 20287 8736
rect 20351 8672 20367 8736
rect 20431 8672 20437 8736
rect 20121 8671 20437 8672
rect 9857 8530 9923 8533
rect 10225 8530 10291 8533
rect 11513 8530 11579 8533
rect 9857 8528 11579 8530
rect 9857 8472 9862 8528
rect 9918 8472 10230 8528
rect 10286 8472 11518 8528
rect 11574 8472 11579 8528
rect 9857 8470 11579 8472
rect 9857 8467 9923 8470
rect 10225 8467 10291 8470
rect 11513 8467 11579 8470
rect 3591 8192 3907 8193
rect 3591 8128 3597 8192
rect 3661 8128 3677 8192
rect 3741 8128 3757 8192
rect 3821 8128 3837 8192
rect 3901 8128 3907 8192
rect 3591 8127 3907 8128
rect 8881 8192 9197 8193
rect 8881 8128 8887 8192
rect 8951 8128 8967 8192
rect 9031 8128 9047 8192
rect 9111 8128 9127 8192
rect 9191 8128 9197 8192
rect 8881 8127 9197 8128
rect 14171 8192 14487 8193
rect 14171 8128 14177 8192
rect 14241 8128 14257 8192
rect 14321 8128 14337 8192
rect 14401 8128 14417 8192
rect 14481 8128 14487 8192
rect 14171 8127 14487 8128
rect 19461 8192 19777 8193
rect 19461 8128 19467 8192
rect 19531 8128 19547 8192
rect 19611 8128 19627 8192
rect 19691 8128 19707 8192
rect 19771 8128 19777 8192
rect 19461 8127 19777 8128
rect 4251 7648 4567 7649
rect 4251 7584 4257 7648
rect 4321 7584 4337 7648
rect 4401 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4567 7648
rect 4251 7583 4567 7584
rect 9541 7648 9857 7649
rect 9541 7584 9547 7648
rect 9611 7584 9627 7648
rect 9691 7584 9707 7648
rect 9771 7584 9787 7648
rect 9851 7584 9857 7648
rect 9541 7583 9857 7584
rect 14831 7648 15147 7649
rect 14831 7584 14837 7648
rect 14901 7584 14917 7648
rect 14981 7584 14997 7648
rect 15061 7584 15077 7648
rect 15141 7584 15147 7648
rect 14831 7583 15147 7584
rect 20121 7648 20437 7649
rect 20121 7584 20127 7648
rect 20191 7584 20207 7648
rect 20271 7584 20287 7648
rect 20351 7584 20367 7648
rect 20431 7584 20437 7648
rect 20121 7583 20437 7584
rect 3591 7104 3907 7105
rect 3591 7040 3597 7104
rect 3661 7040 3677 7104
rect 3741 7040 3757 7104
rect 3821 7040 3837 7104
rect 3901 7040 3907 7104
rect 3591 7039 3907 7040
rect 8881 7104 9197 7105
rect 8881 7040 8887 7104
rect 8951 7040 8967 7104
rect 9031 7040 9047 7104
rect 9111 7040 9127 7104
rect 9191 7040 9197 7104
rect 8881 7039 9197 7040
rect 14171 7104 14487 7105
rect 14171 7040 14177 7104
rect 14241 7040 14257 7104
rect 14321 7040 14337 7104
rect 14401 7040 14417 7104
rect 14481 7040 14487 7104
rect 14171 7039 14487 7040
rect 19461 7104 19777 7105
rect 19461 7040 19467 7104
rect 19531 7040 19547 7104
rect 19611 7040 19627 7104
rect 19691 7040 19707 7104
rect 19771 7040 19777 7104
rect 19461 7039 19777 7040
rect 4251 6560 4567 6561
rect 4251 6496 4257 6560
rect 4321 6496 4337 6560
rect 4401 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4567 6560
rect 4251 6495 4567 6496
rect 9541 6560 9857 6561
rect 9541 6496 9547 6560
rect 9611 6496 9627 6560
rect 9691 6496 9707 6560
rect 9771 6496 9787 6560
rect 9851 6496 9857 6560
rect 9541 6495 9857 6496
rect 14831 6560 15147 6561
rect 14831 6496 14837 6560
rect 14901 6496 14917 6560
rect 14981 6496 14997 6560
rect 15061 6496 15077 6560
rect 15141 6496 15147 6560
rect 14831 6495 15147 6496
rect 20121 6560 20437 6561
rect 20121 6496 20127 6560
rect 20191 6496 20207 6560
rect 20271 6496 20287 6560
rect 20351 6496 20367 6560
rect 20431 6496 20437 6560
rect 20121 6495 20437 6496
rect 3591 6016 3907 6017
rect 3591 5952 3597 6016
rect 3661 5952 3677 6016
rect 3741 5952 3757 6016
rect 3821 5952 3837 6016
rect 3901 5952 3907 6016
rect 3591 5951 3907 5952
rect 8881 6016 9197 6017
rect 8881 5952 8887 6016
rect 8951 5952 8967 6016
rect 9031 5952 9047 6016
rect 9111 5952 9127 6016
rect 9191 5952 9197 6016
rect 8881 5951 9197 5952
rect 14171 6016 14487 6017
rect 14171 5952 14177 6016
rect 14241 5952 14257 6016
rect 14321 5952 14337 6016
rect 14401 5952 14417 6016
rect 14481 5952 14487 6016
rect 14171 5951 14487 5952
rect 19461 6016 19777 6017
rect 19461 5952 19467 6016
rect 19531 5952 19547 6016
rect 19611 5952 19627 6016
rect 19691 5952 19707 6016
rect 19771 5952 19777 6016
rect 19461 5951 19777 5952
rect 9673 5674 9739 5677
rect 11145 5674 11211 5677
rect 9673 5672 11211 5674
rect 9673 5616 9678 5672
rect 9734 5616 11150 5672
rect 11206 5616 11211 5672
rect 9673 5614 11211 5616
rect 9673 5611 9739 5614
rect 11145 5611 11211 5614
rect 4251 5472 4567 5473
rect 4251 5408 4257 5472
rect 4321 5408 4337 5472
rect 4401 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4567 5472
rect 4251 5407 4567 5408
rect 9541 5472 9857 5473
rect 9541 5408 9547 5472
rect 9611 5408 9627 5472
rect 9691 5408 9707 5472
rect 9771 5408 9787 5472
rect 9851 5408 9857 5472
rect 9541 5407 9857 5408
rect 14831 5472 15147 5473
rect 14831 5408 14837 5472
rect 14901 5408 14917 5472
rect 14981 5408 14997 5472
rect 15061 5408 15077 5472
rect 15141 5408 15147 5472
rect 14831 5407 15147 5408
rect 20121 5472 20437 5473
rect 20121 5408 20127 5472
rect 20191 5408 20207 5472
rect 20271 5408 20287 5472
rect 20351 5408 20367 5472
rect 20431 5408 20437 5472
rect 20121 5407 20437 5408
rect 3591 4928 3907 4929
rect 3591 4864 3597 4928
rect 3661 4864 3677 4928
rect 3741 4864 3757 4928
rect 3821 4864 3837 4928
rect 3901 4864 3907 4928
rect 3591 4863 3907 4864
rect 8881 4928 9197 4929
rect 8881 4864 8887 4928
rect 8951 4864 8967 4928
rect 9031 4864 9047 4928
rect 9111 4864 9127 4928
rect 9191 4864 9197 4928
rect 8881 4863 9197 4864
rect 14171 4928 14487 4929
rect 14171 4864 14177 4928
rect 14241 4864 14257 4928
rect 14321 4864 14337 4928
rect 14401 4864 14417 4928
rect 14481 4864 14487 4928
rect 14171 4863 14487 4864
rect 19461 4928 19777 4929
rect 19461 4864 19467 4928
rect 19531 4864 19547 4928
rect 19611 4864 19627 4928
rect 19691 4864 19707 4928
rect 19771 4864 19777 4928
rect 19461 4863 19777 4864
rect 4251 4384 4567 4385
rect 4251 4320 4257 4384
rect 4321 4320 4337 4384
rect 4401 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4567 4384
rect 4251 4319 4567 4320
rect 9541 4384 9857 4385
rect 9541 4320 9547 4384
rect 9611 4320 9627 4384
rect 9691 4320 9707 4384
rect 9771 4320 9787 4384
rect 9851 4320 9857 4384
rect 9541 4319 9857 4320
rect 14831 4384 15147 4385
rect 14831 4320 14837 4384
rect 14901 4320 14917 4384
rect 14981 4320 14997 4384
rect 15061 4320 15077 4384
rect 15141 4320 15147 4384
rect 14831 4319 15147 4320
rect 20121 4384 20437 4385
rect 20121 4320 20127 4384
rect 20191 4320 20207 4384
rect 20271 4320 20287 4384
rect 20351 4320 20367 4384
rect 20431 4320 20437 4384
rect 20121 4319 20437 4320
rect 9765 4178 9831 4181
rect 12985 4178 13051 4181
rect 9765 4176 13051 4178
rect 9765 4120 9770 4176
rect 9826 4120 12990 4176
rect 13046 4120 13051 4176
rect 9765 4118 13051 4120
rect 9765 4115 9831 4118
rect 12985 4115 13051 4118
rect 3591 3840 3907 3841
rect 3591 3776 3597 3840
rect 3661 3776 3677 3840
rect 3741 3776 3757 3840
rect 3821 3776 3837 3840
rect 3901 3776 3907 3840
rect 3591 3775 3907 3776
rect 8881 3840 9197 3841
rect 8881 3776 8887 3840
rect 8951 3776 8967 3840
rect 9031 3776 9047 3840
rect 9111 3776 9127 3840
rect 9191 3776 9197 3840
rect 8881 3775 9197 3776
rect 14171 3840 14487 3841
rect 14171 3776 14177 3840
rect 14241 3776 14257 3840
rect 14321 3776 14337 3840
rect 14401 3776 14417 3840
rect 14481 3776 14487 3840
rect 14171 3775 14487 3776
rect 19461 3840 19777 3841
rect 19461 3776 19467 3840
rect 19531 3776 19547 3840
rect 19611 3776 19627 3840
rect 19691 3776 19707 3840
rect 19771 3776 19777 3840
rect 19461 3775 19777 3776
rect 4251 3296 4567 3297
rect 4251 3232 4257 3296
rect 4321 3232 4337 3296
rect 4401 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4567 3296
rect 4251 3231 4567 3232
rect 9541 3296 9857 3297
rect 9541 3232 9547 3296
rect 9611 3232 9627 3296
rect 9691 3232 9707 3296
rect 9771 3232 9787 3296
rect 9851 3232 9857 3296
rect 9541 3231 9857 3232
rect 14831 3296 15147 3297
rect 14831 3232 14837 3296
rect 14901 3232 14917 3296
rect 14981 3232 14997 3296
rect 15061 3232 15077 3296
rect 15141 3232 15147 3296
rect 14831 3231 15147 3232
rect 20121 3296 20437 3297
rect 20121 3232 20127 3296
rect 20191 3232 20207 3296
rect 20271 3232 20287 3296
rect 20351 3232 20367 3296
rect 20431 3232 20437 3296
rect 20121 3231 20437 3232
rect 3591 2752 3907 2753
rect 3591 2688 3597 2752
rect 3661 2688 3677 2752
rect 3741 2688 3757 2752
rect 3821 2688 3837 2752
rect 3901 2688 3907 2752
rect 3591 2687 3907 2688
rect 8881 2752 9197 2753
rect 8881 2688 8887 2752
rect 8951 2688 8967 2752
rect 9031 2688 9047 2752
rect 9111 2688 9127 2752
rect 9191 2688 9197 2752
rect 8881 2687 9197 2688
rect 14171 2752 14487 2753
rect 14171 2688 14177 2752
rect 14241 2688 14257 2752
rect 14321 2688 14337 2752
rect 14401 2688 14417 2752
rect 14481 2688 14487 2752
rect 14171 2687 14487 2688
rect 19461 2752 19777 2753
rect 19461 2688 19467 2752
rect 19531 2688 19547 2752
rect 19611 2688 19627 2752
rect 19691 2688 19707 2752
rect 19771 2688 19777 2752
rect 19461 2687 19777 2688
rect 4251 2208 4567 2209
rect 4251 2144 4257 2208
rect 4321 2144 4337 2208
rect 4401 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4567 2208
rect 4251 2143 4567 2144
rect 9541 2208 9857 2209
rect 9541 2144 9547 2208
rect 9611 2144 9627 2208
rect 9691 2144 9707 2208
rect 9771 2144 9787 2208
rect 9851 2144 9857 2208
rect 9541 2143 9857 2144
rect 14831 2208 15147 2209
rect 14831 2144 14837 2208
rect 14901 2144 14917 2208
rect 14981 2144 14997 2208
rect 15061 2144 15077 2208
rect 15141 2144 15147 2208
rect 14831 2143 15147 2144
rect 20121 2208 20437 2209
rect 20121 2144 20127 2208
rect 20191 2144 20207 2208
rect 20271 2144 20287 2208
rect 20351 2144 20367 2208
rect 20431 2144 20437 2208
rect 20121 2143 20437 2144
rect 22185 2138 22251 2141
rect 22608 2138 23408 2168
rect 22185 2136 23408 2138
rect 22185 2080 22190 2136
rect 22246 2080 23408 2136
rect 22185 2078 23408 2080
rect 22185 2075 22251 2078
rect 22608 2048 23408 2078
<< via3 >>
rect 4257 22876 4321 22880
rect 4257 22820 4261 22876
rect 4261 22820 4317 22876
rect 4317 22820 4321 22876
rect 4257 22816 4321 22820
rect 4337 22876 4401 22880
rect 4337 22820 4341 22876
rect 4341 22820 4397 22876
rect 4397 22820 4401 22876
rect 4337 22816 4401 22820
rect 4417 22876 4481 22880
rect 4417 22820 4421 22876
rect 4421 22820 4477 22876
rect 4477 22820 4481 22876
rect 4417 22816 4481 22820
rect 4497 22876 4561 22880
rect 4497 22820 4501 22876
rect 4501 22820 4557 22876
rect 4557 22820 4561 22876
rect 4497 22816 4561 22820
rect 9547 22876 9611 22880
rect 9547 22820 9551 22876
rect 9551 22820 9607 22876
rect 9607 22820 9611 22876
rect 9547 22816 9611 22820
rect 9627 22876 9691 22880
rect 9627 22820 9631 22876
rect 9631 22820 9687 22876
rect 9687 22820 9691 22876
rect 9627 22816 9691 22820
rect 9707 22876 9771 22880
rect 9707 22820 9711 22876
rect 9711 22820 9767 22876
rect 9767 22820 9771 22876
rect 9707 22816 9771 22820
rect 9787 22876 9851 22880
rect 9787 22820 9791 22876
rect 9791 22820 9847 22876
rect 9847 22820 9851 22876
rect 9787 22816 9851 22820
rect 14837 22876 14901 22880
rect 14837 22820 14841 22876
rect 14841 22820 14897 22876
rect 14897 22820 14901 22876
rect 14837 22816 14901 22820
rect 14917 22876 14981 22880
rect 14917 22820 14921 22876
rect 14921 22820 14977 22876
rect 14977 22820 14981 22876
rect 14917 22816 14981 22820
rect 14997 22876 15061 22880
rect 14997 22820 15001 22876
rect 15001 22820 15057 22876
rect 15057 22820 15061 22876
rect 14997 22816 15061 22820
rect 15077 22876 15141 22880
rect 15077 22820 15081 22876
rect 15081 22820 15137 22876
rect 15137 22820 15141 22876
rect 15077 22816 15141 22820
rect 20127 22876 20191 22880
rect 20127 22820 20131 22876
rect 20131 22820 20187 22876
rect 20187 22820 20191 22876
rect 20127 22816 20191 22820
rect 20207 22876 20271 22880
rect 20207 22820 20211 22876
rect 20211 22820 20267 22876
rect 20267 22820 20271 22876
rect 20207 22816 20271 22820
rect 20287 22876 20351 22880
rect 20287 22820 20291 22876
rect 20291 22820 20347 22876
rect 20347 22820 20351 22876
rect 20287 22816 20351 22820
rect 20367 22876 20431 22880
rect 20367 22820 20371 22876
rect 20371 22820 20427 22876
rect 20427 22820 20431 22876
rect 20367 22816 20431 22820
rect 3597 22332 3661 22336
rect 3597 22276 3601 22332
rect 3601 22276 3657 22332
rect 3657 22276 3661 22332
rect 3597 22272 3661 22276
rect 3677 22332 3741 22336
rect 3677 22276 3681 22332
rect 3681 22276 3737 22332
rect 3737 22276 3741 22332
rect 3677 22272 3741 22276
rect 3757 22332 3821 22336
rect 3757 22276 3761 22332
rect 3761 22276 3817 22332
rect 3817 22276 3821 22332
rect 3757 22272 3821 22276
rect 3837 22332 3901 22336
rect 3837 22276 3841 22332
rect 3841 22276 3897 22332
rect 3897 22276 3901 22332
rect 3837 22272 3901 22276
rect 8887 22332 8951 22336
rect 8887 22276 8891 22332
rect 8891 22276 8947 22332
rect 8947 22276 8951 22332
rect 8887 22272 8951 22276
rect 8967 22332 9031 22336
rect 8967 22276 8971 22332
rect 8971 22276 9027 22332
rect 9027 22276 9031 22332
rect 8967 22272 9031 22276
rect 9047 22332 9111 22336
rect 9047 22276 9051 22332
rect 9051 22276 9107 22332
rect 9107 22276 9111 22332
rect 9047 22272 9111 22276
rect 9127 22332 9191 22336
rect 9127 22276 9131 22332
rect 9131 22276 9187 22332
rect 9187 22276 9191 22332
rect 9127 22272 9191 22276
rect 14177 22332 14241 22336
rect 14177 22276 14181 22332
rect 14181 22276 14237 22332
rect 14237 22276 14241 22332
rect 14177 22272 14241 22276
rect 14257 22332 14321 22336
rect 14257 22276 14261 22332
rect 14261 22276 14317 22332
rect 14317 22276 14321 22332
rect 14257 22272 14321 22276
rect 14337 22332 14401 22336
rect 14337 22276 14341 22332
rect 14341 22276 14397 22332
rect 14397 22276 14401 22332
rect 14337 22272 14401 22276
rect 14417 22332 14481 22336
rect 14417 22276 14421 22332
rect 14421 22276 14477 22332
rect 14477 22276 14481 22332
rect 14417 22272 14481 22276
rect 19467 22332 19531 22336
rect 19467 22276 19471 22332
rect 19471 22276 19527 22332
rect 19527 22276 19531 22332
rect 19467 22272 19531 22276
rect 19547 22332 19611 22336
rect 19547 22276 19551 22332
rect 19551 22276 19607 22332
rect 19607 22276 19611 22332
rect 19547 22272 19611 22276
rect 19627 22332 19691 22336
rect 19627 22276 19631 22332
rect 19631 22276 19687 22332
rect 19687 22276 19691 22332
rect 19627 22272 19691 22276
rect 19707 22332 19771 22336
rect 19707 22276 19711 22332
rect 19711 22276 19767 22332
rect 19767 22276 19771 22332
rect 19707 22272 19771 22276
rect 4257 21788 4321 21792
rect 4257 21732 4261 21788
rect 4261 21732 4317 21788
rect 4317 21732 4321 21788
rect 4257 21728 4321 21732
rect 4337 21788 4401 21792
rect 4337 21732 4341 21788
rect 4341 21732 4397 21788
rect 4397 21732 4401 21788
rect 4337 21728 4401 21732
rect 4417 21788 4481 21792
rect 4417 21732 4421 21788
rect 4421 21732 4477 21788
rect 4477 21732 4481 21788
rect 4417 21728 4481 21732
rect 4497 21788 4561 21792
rect 4497 21732 4501 21788
rect 4501 21732 4557 21788
rect 4557 21732 4561 21788
rect 4497 21728 4561 21732
rect 9547 21788 9611 21792
rect 9547 21732 9551 21788
rect 9551 21732 9607 21788
rect 9607 21732 9611 21788
rect 9547 21728 9611 21732
rect 9627 21788 9691 21792
rect 9627 21732 9631 21788
rect 9631 21732 9687 21788
rect 9687 21732 9691 21788
rect 9627 21728 9691 21732
rect 9707 21788 9771 21792
rect 9707 21732 9711 21788
rect 9711 21732 9767 21788
rect 9767 21732 9771 21788
rect 9707 21728 9771 21732
rect 9787 21788 9851 21792
rect 9787 21732 9791 21788
rect 9791 21732 9847 21788
rect 9847 21732 9851 21788
rect 9787 21728 9851 21732
rect 14837 21788 14901 21792
rect 14837 21732 14841 21788
rect 14841 21732 14897 21788
rect 14897 21732 14901 21788
rect 14837 21728 14901 21732
rect 14917 21788 14981 21792
rect 14917 21732 14921 21788
rect 14921 21732 14977 21788
rect 14977 21732 14981 21788
rect 14917 21728 14981 21732
rect 14997 21788 15061 21792
rect 14997 21732 15001 21788
rect 15001 21732 15057 21788
rect 15057 21732 15061 21788
rect 14997 21728 15061 21732
rect 15077 21788 15141 21792
rect 15077 21732 15081 21788
rect 15081 21732 15137 21788
rect 15137 21732 15141 21788
rect 15077 21728 15141 21732
rect 20127 21788 20191 21792
rect 20127 21732 20131 21788
rect 20131 21732 20187 21788
rect 20187 21732 20191 21788
rect 20127 21728 20191 21732
rect 20207 21788 20271 21792
rect 20207 21732 20211 21788
rect 20211 21732 20267 21788
rect 20267 21732 20271 21788
rect 20207 21728 20271 21732
rect 20287 21788 20351 21792
rect 20287 21732 20291 21788
rect 20291 21732 20347 21788
rect 20347 21732 20351 21788
rect 20287 21728 20351 21732
rect 20367 21788 20431 21792
rect 20367 21732 20371 21788
rect 20371 21732 20427 21788
rect 20427 21732 20431 21788
rect 20367 21728 20431 21732
rect 3597 21244 3661 21248
rect 3597 21188 3601 21244
rect 3601 21188 3657 21244
rect 3657 21188 3661 21244
rect 3597 21184 3661 21188
rect 3677 21244 3741 21248
rect 3677 21188 3681 21244
rect 3681 21188 3737 21244
rect 3737 21188 3741 21244
rect 3677 21184 3741 21188
rect 3757 21244 3821 21248
rect 3757 21188 3761 21244
rect 3761 21188 3817 21244
rect 3817 21188 3821 21244
rect 3757 21184 3821 21188
rect 3837 21244 3901 21248
rect 3837 21188 3841 21244
rect 3841 21188 3897 21244
rect 3897 21188 3901 21244
rect 3837 21184 3901 21188
rect 8887 21244 8951 21248
rect 8887 21188 8891 21244
rect 8891 21188 8947 21244
rect 8947 21188 8951 21244
rect 8887 21184 8951 21188
rect 8967 21244 9031 21248
rect 8967 21188 8971 21244
rect 8971 21188 9027 21244
rect 9027 21188 9031 21244
rect 8967 21184 9031 21188
rect 9047 21244 9111 21248
rect 9047 21188 9051 21244
rect 9051 21188 9107 21244
rect 9107 21188 9111 21244
rect 9047 21184 9111 21188
rect 9127 21244 9191 21248
rect 9127 21188 9131 21244
rect 9131 21188 9187 21244
rect 9187 21188 9191 21244
rect 9127 21184 9191 21188
rect 14177 21244 14241 21248
rect 14177 21188 14181 21244
rect 14181 21188 14237 21244
rect 14237 21188 14241 21244
rect 14177 21184 14241 21188
rect 14257 21244 14321 21248
rect 14257 21188 14261 21244
rect 14261 21188 14317 21244
rect 14317 21188 14321 21244
rect 14257 21184 14321 21188
rect 14337 21244 14401 21248
rect 14337 21188 14341 21244
rect 14341 21188 14397 21244
rect 14397 21188 14401 21244
rect 14337 21184 14401 21188
rect 14417 21244 14481 21248
rect 14417 21188 14421 21244
rect 14421 21188 14477 21244
rect 14477 21188 14481 21244
rect 14417 21184 14481 21188
rect 19467 21244 19531 21248
rect 19467 21188 19471 21244
rect 19471 21188 19527 21244
rect 19527 21188 19531 21244
rect 19467 21184 19531 21188
rect 19547 21244 19611 21248
rect 19547 21188 19551 21244
rect 19551 21188 19607 21244
rect 19607 21188 19611 21244
rect 19547 21184 19611 21188
rect 19627 21244 19691 21248
rect 19627 21188 19631 21244
rect 19631 21188 19687 21244
rect 19687 21188 19691 21244
rect 19627 21184 19691 21188
rect 19707 21244 19771 21248
rect 19707 21188 19711 21244
rect 19711 21188 19767 21244
rect 19767 21188 19771 21244
rect 19707 21184 19771 21188
rect 4257 20700 4321 20704
rect 4257 20644 4261 20700
rect 4261 20644 4317 20700
rect 4317 20644 4321 20700
rect 4257 20640 4321 20644
rect 4337 20700 4401 20704
rect 4337 20644 4341 20700
rect 4341 20644 4397 20700
rect 4397 20644 4401 20700
rect 4337 20640 4401 20644
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 9547 20700 9611 20704
rect 9547 20644 9551 20700
rect 9551 20644 9607 20700
rect 9607 20644 9611 20700
rect 9547 20640 9611 20644
rect 9627 20700 9691 20704
rect 9627 20644 9631 20700
rect 9631 20644 9687 20700
rect 9687 20644 9691 20700
rect 9627 20640 9691 20644
rect 9707 20700 9771 20704
rect 9707 20644 9711 20700
rect 9711 20644 9767 20700
rect 9767 20644 9771 20700
rect 9707 20640 9771 20644
rect 9787 20700 9851 20704
rect 9787 20644 9791 20700
rect 9791 20644 9847 20700
rect 9847 20644 9851 20700
rect 9787 20640 9851 20644
rect 14837 20700 14901 20704
rect 14837 20644 14841 20700
rect 14841 20644 14897 20700
rect 14897 20644 14901 20700
rect 14837 20640 14901 20644
rect 14917 20700 14981 20704
rect 14917 20644 14921 20700
rect 14921 20644 14977 20700
rect 14977 20644 14981 20700
rect 14917 20640 14981 20644
rect 14997 20700 15061 20704
rect 14997 20644 15001 20700
rect 15001 20644 15057 20700
rect 15057 20644 15061 20700
rect 14997 20640 15061 20644
rect 15077 20700 15141 20704
rect 15077 20644 15081 20700
rect 15081 20644 15137 20700
rect 15137 20644 15141 20700
rect 15077 20640 15141 20644
rect 20127 20700 20191 20704
rect 20127 20644 20131 20700
rect 20131 20644 20187 20700
rect 20187 20644 20191 20700
rect 20127 20640 20191 20644
rect 20207 20700 20271 20704
rect 20207 20644 20211 20700
rect 20211 20644 20267 20700
rect 20267 20644 20271 20700
rect 20207 20640 20271 20644
rect 20287 20700 20351 20704
rect 20287 20644 20291 20700
rect 20291 20644 20347 20700
rect 20347 20644 20351 20700
rect 20287 20640 20351 20644
rect 20367 20700 20431 20704
rect 20367 20644 20371 20700
rect 20371 20644 20427 20700
rect 20427 20644 20431 20700
rect 20367 20640 20431 20644
rect 3597 20156 3661 20160
rect 3597 20100 3601 20156
rect 3601 20100 3657 20156
rect 3657 20100 3661 20156
rect 3597 20096 3661 20100
rect 3677 20156 3741 20160
rect 3677 20100 3681 20156
rect 3681 20100 3737 20156
rect 3737 20100 3741 20156
rect 3677 20096 3741 20100
rect 3757 20156 3821 20160
rect 3757 20100 3761 20156
rect 3761 20100 3817 20156
rect 3817 20100 3821 20156
rect 3757 20096 3821 20100
rect 3837 20156 3901 20160
rect 3837 20100 3841 20156
rect 3841 20100 3897 20156
rect 3897 20100 3901 20156
rect 3837 20096 3901 20100
rect 8887 20156 8951 20160
rect 8887 20100 8891 20156
rect 8891 20100 8947 20156
rect 8947 20100 8951 20156
rect 8887 20096 8951 20100
rect 8967 20156 9031 20160
rect 8967 20100 8971 20156
rect 8971 20100 9027 20156
rect 9027 20100 9031 20156
rect 8967 20096 9031 20100
rect 9047 20156 9111 20160
rect 9047 20100 9051 20156
rect 9051 20100 9107 20156
rect 9107 20100 9111 20156
rect 9047 20096 9111 20100
rect 9127 20156 9191 20160
rect 9127 20100 9131 20156
rect 9131 20100 9187 20156
rect 9187 20100 9191 20156
rect 9127 20096 9191 20100
rect 14177 20156 14241 20160
rect 14177 20100 14181 20156
rect 14181 20100 14237 20156
rect 14237 20100 14241 20156
rect 14177 20096 14241 20100
rect 14257 20156 14321 20160
rect 14257 20100 14261 20156
rect 14261 20100 14317 20156
rect 14317 20100 14321 20156
rect 14257 20096 14321 20100
rect 14337 20156 14401 20160
rect 14337 20100 14341 20156
rect 14341 20100 14397 20156
rect 14397 20100 14401 20156
rect 14337 20096 14401 20100
rect 14417 20156 14481 20160
rect 14417 20100 14421 20156
rect 14421 20100 14477 20156
rect 14477 20100 14481 20156
rect 14417 20096 14481 20100
rect 19467 20156 19531 20160
rect 19467 20100 19471 20156
rect 19471 20100 19527 20156
rect 19527 20100 19531 20156
rect 19467 20096 19531 20100
rect 19547 20156 19611 20160
rect 19547 20100 19551 20156
rect 19551 20100 19607 20156
rect 19607 20100 19611 20156
rect 19547 20096 19611 20100
rect 19627 20156 19691 20160
rect 19627 20100 19631 20156
rect 19631 20100 19687 20156
rect 19687 20100 19691 20156
rect 19627 20096 19691 20100
rect 19707 20156 19771 20160
rect 19707 20100 19711 20156
rect 19711 20100 19767 20156
rect 19767 20100 19771 20156
rect 19707 20096 19771 20100
rect 4257 19612 4321 19616
rect 4257 19556 4261 19612
rect 4261 19556 4317 19612
rect 4317 19556 4321 19612
rect 4257 19552 4321 19556
rect 4337 19612 4401 19616
rect 4337 19556 4341 19612
rect 4341 19556 4397 19612
rect 4397 19556 4401 19612
rect 4337 19552 4401 19556
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 9547 19612 9611 19616
rect 9547 19556 9551 19612
rect 9551 19556 9607 19612
rect 9607 19556 9611 19612
rect 9547 19552 9611 19556
rect 9627 19612 9691 19616
rect 9627 19556 9631 19612
rect 9631 19556 9687 19612
rect 9687 19556 9691 19612
rect 9627 19552 9691 19556
rect 9707 19612 9771 19616
rect 9707 19556 9711 19612
rect 9711 19556 9767 19612
rect 9767 19556 9771 19612
rect 9707 19552 9771 19556
rect 9787 19612 9851 19616
rect 9787 19556 9791 19612
rect 9791 19556 9847 19612
rect 9847 19556 9851 19612
rect 9787 19552 9851 19556
rect 14837 19612 14901 19616
rect 14837 19556 14841 19612
rect 14841 19556 14897 19612
rect 14897 19556 14901 19612
rect 14837 19552 14901 19556
rect 14917 19612 14981 19616
rect 14917 19556 14921 19612
rect 14921 19556 14977 19612
rect 14977 19556 14981 19612
rect 14917 19552 14981 19556
rect 14997 19612 15061 19616
rect 14997 19556 15001 19612
rect 15001 19556 15057 19612
rect 15057 19556 15061 19612
rect 14997 19552 15061 19556
rect 15077 19612 15141 19616
rect 15077 19556 15081 19612
rect 15081 19556 15137 19612
rect 15137 19556 15141 19612
rect 15077 19552 15141 19556
rect 20127 19612 20191 19616
rect 20127 19556 20131 19612
rect 20131 19556 20187 19612
rect 20187 19556 20191 19612
rect 20127 19552 20191 19556
rect 20207 19612 20271 19616
rect 20207 19556 20211 19612
rect 20211 19556 20267 19612
rect 20267 19556 20271 19612
rect 20207 19552 20271 19556
rect 20287 19612 20351 19616
rect 20287 19556 20291 19612
rect 20291 19556 20347 19612
rect 20347 19556 20351 19612
rect 20287 19552 20351 19556
rect 20367 19612 20431 19616
rect 20367 19556 20371 19612
rect 20371 19556 20427 19612
rect 20427 19556 20431 19612
rect 20367 19552 20431 19556
rect 3597 19068 3661 19072
rect 3597 19012 3601 19068
rect 3601 19012 3657 19068
rect 3657 19012 3661 19068
rect 3597 19008 3661 19012
rect 3677 19068 3741 19072
rect 3677 19012 3681 19068
rect 3681 19012 3737 19068
rect 3737 19012 3741 19068
rect 3677 19008 3741 19012
rect 3757 19068 3821 19072
rect 3757 19012 3761 19068
rect 3761 19012 3817 19068
rect 3817 19012 3821 19068
rect 3757 19008 3821 19012
rect 3837 19068 3901 19072
rect 3837 19012 3841 19068
rect 3841 19012 3897 19068
rect 3897 19012 3901 19068
rect 3837 19008 3901 19012
rect 8887 19068 8951 19072
rect 8887 19012 8891 19068
rect 8891 19012 8947 19068
rect 8947 19012 8951 19068
rect 8887 19008 8951 19012
rect 8967 19068 9031 19072
rect 8967 19012 8971 19068
rect 8971 19012 9027 19068
rect 9027 19012 9031 19068
rect 8967 19008 9031 19012
rect 9047 19068 9111 19072
rect 9047 19012 9051 19068
rect 9051 19012 9107 19068
rect 9107 19012 9111 19068
rect 9047 19008 9111 19012
rect 9127 19068 9191 19072
rect 9127 19012 9131 19068
rect 9131 19012 9187 19068
rect 9187 19012 9191 19068
rect 9127 19008 9191 19012
rect 14177 19068 14241 19072
rect 14177 19012 14181 19068
rect 14181 19012 14237 19068
rect 14237 19012 14241 19068
rect 14177 19008 14241 19012
rect 14257 19068 14321 19072
rect 14257 19012 14261 19068
rect 14261 19012 14317 19068
rect 14317 19012 14321 19068
rect 14257 19008 14321 19012
rect 14337 19068 14401 19072
rect 14337 19012 14341 19068
rect 14341 19012 14397 19068
rect 14397 19012 14401 19068
rect 14337 19008 14401 19012
rect 14417 19068 14481 19072
rect 14417 19012 14421 19068
rect 14421 19012 14477 19068
rect 14477 19012 14481 19068
rect 14417 19008 14481 19012
rect 19467 19068 19531 19072
rect 19467 19012 19471 19068
rect 19471 19012 19527 19068
rect 19527 19012 19531 19068
rect 19467 19008 19531 19012
rect 19547 19068 19611 19072
rect 19547 19012 19551 19068
rect 19551 19012 19607 19068
rect 19607 19012 19611 19068
rect 19547 19008 19611 19012
rect 19627 19068 19691 19072
rect 19627 19012 19631 19068
rect 19631 19012 19687 19068
rect 19687 19012 19691 19068
rect 19627 19008 19691 19012
rect 19707 19068 19771 19072
rect 19707 19012 19711 19068
rect 19711 19012 19767 19068
rect 19767 19012 19771 19068
rect 19707 19008 19771 19012
rect 4257 18524 4321 18528
rect 4257 18468 4261 18524
rect 4261 18468 4317 18524
rect 4317 18468 4321 18524
rect 4257 18464 4321 18468
rect 4337 18524 4401 18528
rect 4337 18468 4341 18524
rect 4341 18468 4397 18524
rect 4397 18468 4401 18524
rect 4337 18464 4401 18468
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 9547 18524 9611 18528
rect 9547 18468 9551 18524
rect 9551 18468 9607 18524
rect 9607 18468 9611 18524
rect 9547 18464 9611 18468
rect 9627 18524 9691 18528
rect 9627 18468 9631 18524
rect 9631 18468 9687 18524
rect 9687 18468 9691 18524
rect 9627 18464 9691 18468
rect 9707 18524 9771 18528
rect 9707 18468 9711 18524
rect 9711 18468 9767 18524
rect 9767 18468 9771 18524
rect 9707 18464 9771 18468
rect 9787 18524 9851 18528
rect 9787 18468 9791 18524
rect 9791 18468 9847 18524
rect 9847 18468 9851 18524
rect 9787 18464 9851 18468
rect 14837 18524 14901 18528
rect 14837 18468 14841 18524
rect 14841 18468 14897 18524
rect 14897 18468 14901 18524
rect 14837 18464 14901 18468
rect 14917 18524 14981 18528
rect 14917 18468 14921 18524
rect 14921 18468 14977 18524
rect 14977 18468 14981 18524
rect 14917 18464 14981 18468
rect 14997 18524 15061 18528
rect 14997 18468 15001 18524
rect 15001 18468 15057 18524
rect 15057 18468 15061 18524
rect 14997 18464 15061 18468
rect 15077 18524 15141 18528
rect 15077 18468 15081 18524
rect 15081 18468 15137 18524
rect 15137 18468 15141 18524
rect 15077 18464 15141 18468
rect 20127 18524 20191 18528
rect 20127 18468 20131 18524
rect 20131 18468 20187 18524
rect 20187 18468 20191 18524
rect 20127 18464 20191 18468
rect 20207 18524 20271 18528
rect 20207 18468 20211 18524
rect 20211 18468 20267 18524
rect 20267 18468 20271 18524
rect 20207 18464 20271 18468
rect 20287 18524 20351 18528
rect 20287 18468 20291 18524
rect 20291 18468 20347 18524
rect 20347 18468 20351 18524
rect 20287 18464 20351 18468
rect 20367 18524 20431 18528
rect 20367 18468 20371 18524
rect 20371 18468 20427 18524
rect 20427 18468 20431 18524
rect 20367 18464 20431 18468
rect 3597 17980 3661 17984
rect 3597 17924 3601 17980
rect 3601 17924 3657 17980
rect 3657 17924 3661 17980
rect 3597 17920 3661 17924
rect 3677 17980 3741 17984
rect 3677 17924 3681 17980
rect 3681 17924 3737 17980
rect 3737 17924 3741 17980
rect 3677 17920 3741 17924
rect 3757 17980 3821 17984
rect 3757 17924 3761 17980
rect 3761 17924 3817 17980
rect 3817 17924 3821 17980
rect 3757 17920 3821 17924
rect 3837 17980 3901 17984
rect 3837 17924 3841 17980
rect 3841 17924 3897 17980
rect 3897 17924 3901 17980
rect 3837 17920 3901 17924
rect 8887 17980 8951 17984
rect 8887 17924 8891 17980
rect 8891 17924 8947 17980
rect 8947 17924 8951 17980
rect 8887 17920 8951 17924
rect 8967 17980 9031 17984
rect 8967 17924 8971 17980
rect 8971 17924 9027 17980
rect 9027 17924 9031 17980
rect 8967 17920 9031 17924
rect 9047 17980 9111 17984
rect 9047 17924 9051 17980
rect 9051 17924 9107 17980
rect 9107 17924 9111 17980
rect 9047 17920 9111 17924
rect 9127 17980 9191 17984
rect 9127 17924 9131 17980
rect 9131 17924 9187 17980
rect 9187 17924 9191 17980
rect 9127 17920 9191 17924
rect 14177 17980 14241 17984
rect 14177 17924 14181 17980
rect 14181 17924 14237 17980
rect 14237 17924 14241 17980
rect 14177 17920 14241 17924
rect 14257 17980 14321 17984
rect 14257 17924 14261 17980
rect 14261 17924 14317 17980
rect 14317 17924 14321 17980
rect 14257 17920 14321 17924
rect 14337 17980 14401 17984
rect 14337 17924 14341 17980
rect 14341 17924 14397 17980
rect 14397 17924 14401 17980
rect 14337 17920 14401 17924
rect 14417 17980 14481 17984
rect 14417 17924 14421 17980
rect 14421 17924 14477 17980
rect 14477 17924 14481 17980
rect 14417 17920 14481 17924
rect 19467 17980 19531 17984
rect 19467 17924 19471 17980
rect 19471 17924 19527 17980
rect 19527 17924 19531 17980
rect 19467 17920 19531 17924
rect 19547 17980 19611 17984
rect 19547 17924 19551 17980
rect 19551 17924 19607 17980
rect 19607 17924 19611 17980
rect 19547 17920 19611 17924
rect 19627 17980 19691 17984
rect 19627 17924 19631 17980
rect 19631 17924 19687 17980
rect 19687 17924 19691 17980
rect 19627 17920 19691 17924
rect 19707 17980 19771 17984
rect 19707 17924 19711 17980
rect 19711 17924 19767 17980
rect 19767 17924 19771 17980
rect 19707 17920 19771 17924
rect 4257 17436 4321 17440
rect 4257 17380 4261 17436
rect 4261 17380 4317 17436
rect 4317 17380 4321 17436
rect 4257 17376 4321 17380
rect 4337 17436 4401 17440
rect 4337 17380 4341 17436
rect 4341 17380 4397 17436
rect 4397 17380 4401 17436
rect 4337 17376 4401 17380
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 9547 17436 9611 17440
rect 9547 17380 9551 17436
rect 9551 17380 9607 17436
rect 9607 17380 9611 17436
rect 9547 17376 9611 17380
rect 9627 17436 9691 17440
rect 9627 17380 9631 17436
rect 9631 17380 9687 17436
rect 9687 17380 9691 17436
rect 9627 17376 9691 17380
rect 9707 17436 9771 17440
rect 9707 17380 9711 17436
rect 9711 17380 9767 17436
rect 9767 17380 9771 17436
rect 9707 17376 9771 17380
rect 9787 17436 9851 17440
rect 9787 17380 9791 17436
rect 9791 17380 9847 17436
rect 9847 17380 9851 17436
rect 9787 17376 9851 17380
rect 14837 17436 14901 17440
rect 14837 17380 14841 17436
rect 14841 17380 14897 17436
rect 14897 17380 14901 17436
rect 14837 17376 14901 17380
rect 14917 17436 14981 17440
rect 14917 17380 14921 17436
rect 14921 17380 14977 17436
rect 14977 17380 14981 17436
rect 14917 17376 14981 17380
rect 14997 17436 15061 17440
rect 14997 17380 15001 17436
rect 15001 17380 15057 17436
rect 15057 17380 15061 17436
rect 14997 17376 15061 17380
rect 15077 17436 15141 17440
rect 15077 17380 15081 17436
rect 15081 17380 15137 17436
rect 15137 17380 15141 17436
rect 15077 17376 15141 17380
rect 20127 17436 20191 17440
rect 20127 17380 20131 17436
rect 20131 17380 20187 17436
rect 20187 17380 20191 17436
rect 20127 17376 20191 17380
rect 20207 17436 20271 17440
rect 20207 17380 20211 17436
rect 20211 17380 20267 17436
rect 20267 17380 20271 17436
rect 20207 17376 20271 17380
rect 20287 17436 20351 17440
rect 20287 17380 20291 17436
rect 20291 17380 20347 17436
rect 20347 17380 20351 17436
rect 20287 17376 20351 17380
rect 20367 17436 20431 17440
rect 20367 17380 20371 17436
rect 20371 17380 20427 17436
rect 20427 17380 20431 17436
rect 20367 17376 20431 17380
rect 3597 16892 3661 16896
rect 3597 16836 3601 16892
rect 3601 16836 3657 16892
rect 3657 16836 3661 16892
rect 3597 16832 3661 16836
rect 3677 16892 3741 16896
rect 3677 16836 3681 16892
rect 3681 16836 3737 16892
rect 3737 16836 3741 16892
rect 3677 16832 3741 16836
rect 3757 16892 3821 16896
rect 3757 16836 3761 16892
rect 3761 16836 3817 16892
rect 3817 16836 3821 16892
rect 3757 16832 3821 16836
rect 3837 16892 3901 16896
rect 3837 16836 3841 16892
rect 3841 16836 3897 16892
rect 3897 16836 3901 16892
rect 3837 16832 3901 16836
rect 8887 16892 8951 16896
rect 8887 16836 8891 16892
rect 8891 16836 8947 16892
rect 8947 16836 8951 16892
rect 8887 16832 8951 16836
rect 8967 16892 9031 16896
rect 8967 16836 8971 16892
rect 8971 16836 9027 16892
rect 9027 16836 9031 16892
rect 8967 16832 9031 16836
rect 9047 16892 9111 16896
rect 9047 16836 9051 16892
rect 9051 16836 9107 16892
rect 9107 16836 9111 16892
rect 9047 16832 9111 16836
rect 9127 16892 9191 16896
rect 9127 16836 9131 16892
rect 9131 16836 9187 16892
rect 9187 16836 9191 16892
rect 9127 16832 9191 16836
rect 14177 16892 14241 16896
rect 14177 16836 14181 16892
rect 14181 16836 14237 16892
rect 14237 16836 14241 16892
rect 14177 16832 14241 16836
rect 14257 16892 14321 16896
rect 14257 16836 14261 16892
rect 14261 16836 14317 16892
rect 14317 16836 14321 16892
rect 14257 16832 14321 16836
rect 14337 16892 14401 16896
rect 14337 16836 14341 16892
rect 14341 16836 14397 16892
rect 14397 16836 14401 16892
rect 14337 16832 14401 16836
rect 14417 16892 14481 16896
rect 14417 16836 14421 16892
rect 14421 16836 14477 16892
rect 14477 16836 14481 16892
rect 14417 16832 14481 16836
rect 19467 16892 19531 16896
rect 19467 16836 19471 16892
rect 19471 16836 19527 16892
rect 19527 16836 19531 16892
rect 19467 16832 19531 16836
rect 19547 16892 19611 16896
rect 19547 16836 19551 16892
rect 19551 16836 19607 16892
rect 19607 16836 19611 16892
rect 19547 16832 19611 16836
rect 19627 16892 19691 16896
rect 19627 16836 19631 16892
rect 19631 16836 19687 16892
rect 19687 16836 19691 16892
rect 19627 16832 19691 16836
rect 19707 16892 19771 16896
rect 19707 16836 19711 16892
rect 19711 16836 19767 16892
rect 19767 16836 19771 16892
rect 19707 16832 19771 16836
rect 4257 16348 4321 16352
rect 4257 16292 4261 16348
rect 4261 16292 4317 16348
rect 4317 16292 4321 16348
rect 4257 16288 4321 16292
rect 4337 16348 4401 16352
rect 4337 16292 4341 16348
rect 4341 16292 4397 16348
rect 4397 16292 4401 16348
rect 4337 16288 4401 16292
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 9547 16348 9611 16352
rect 9547 16292 9551 16348
rect 9551 16292 9607 16348
rect 9607 16292 9611 16348
rect 9547 16288 9611 16292
rect 9627 16348 9691 16352
rect 9627 16292 9631 16348
rect 9631 16292 9687 16348
rect 9687 16292 9691 16348
rect 9627 16288 9691 16292
rect 9707 16348 9771 16352
rect 9707 16292 9711 16348
rect 9711 16292 9767 16348
rect 9767 16292 9771 16348
rect 9707 16288 9771 16292
rect 9787 16348 9851 16352
rect 9787 16292 9791 16348
rect 9791 16292 9847 16348
rect 9847 16292 9851 16348
rect 9787 16288 9851 16292
rect 14837 16348 14901 16352
rect 14837 16292 14841 16348
rect 14841 16292 14897 16348
rect 14897 16292 14901 16348
rect 14837 16288 14901 16292
rect 14917 16348 14981 16352
rect 14917 16292 14921 16348
rect 14921 16292 14977 16348
rect 14977 16292 14981 16348
rect 14917 16288 14981 16292
rect 14997 16348 15061 16352
rect 14997 16292 15001 16348
rect 15001 16292 15057 16348
rect 15057 16292 15061 16348
rect 14997 16288 15061 16292
rect 15077 16348 15141 16352
rect 15077 16292 15081 16348
rect 15081 16292 15137 16348
rect 15137 16292 15141 16348
rect 15077 16288 15141 16292
rect 20127 16348 20191 16352
rect 20127 16292 20131 16348
rect 20131 16292 20187 16348
rect 20187 16292 20191 16348
rect 20127 16288 20191 16292
rect 20207 16348 20271 16352
rect 20207 16292 20211 16348
rect 20211 16292 20267 16348
rect 20267 16292 20271 16348
rect 20207 16288 20271 16292
rect 20287 16348 20351 16352
rect 20287 16292 20291 16348
rect 20291 16292 20347 16348
rect 20347 16292 20351 16348
rect 20287 16288 20351 16292
rect 20367 16348 20431 16352
rect 20367 16292 20371 16348
rect 20371 16292 20427 16348
rect 20427 16292 20431 16348
rect 20367 16288 20431 16292
rect 3597 15804 3661 15808
rect 3597 15748 3601 15804
rect 3601 15748 3657 15804
rect 3657 15748 3661 15804
rect 3597 15744 3661 15748
rect 3677 15804 3741 15808
rect 3677 15748 3681 15804
rect 3681 15748 3737 15804
rect 3737 15748 3741 15804
rect 3677 15744 3741 15748
rect 3757 15804 3821 15808
rect 3757 15748 3761 15804
rect 3761 15748 3817 15804
rect 3817 15748 3821 15804
rect 3757 15744 3821 15748
rect 3837 15804 3901 15808
rect 3837 15748 3841 15804
rect 3841 15748 3897 15804
rect 3897 15748 3901 15804
rect 3837 15744 3901 15748
rect 8887 15804 8951 15808
rect 8887 15748 8891 15804
rect 8891 15748 8947 15804
rect 8947 15748 8951 15804
rect 8887 15744 8951 15748
rect 8967 15804 9031 15808
rect 8967 15748 8971 15804
rect 8971 15748 9027 15804
rect 9027 15748 9031 15804
rect 8967 15744 9031 15748
rect 9047 15804 9111 15808
rect 9047 15748 9051 15804
rect 9051 15748 9107 15804
rect 9107 15748 9111 15804
rect 9047 15744 9111 15748
rect 9127 15804 9191 15808
rect 9127 15748 9131 15804
rect 9131 15748 9187 15804
rect 9187 15748 9191 15804
rect 9127 15744 9191 15748
rect 14177 15804 14241 15808
rect 14177 15748 14181 15804
rect 14181 15748 14237 15804
rect 14237 15748 14241 15804
rect 14177 15744 14241 15748
rect 14257 15804 14321 15808
rect 14257 15748 14261 15804
rect 14261 15748 14317 15804
rect 14317 15748 14321 15804
rect 14257 15744 14321 15748
rect 14337 15804 14401 15808
rect 14337 15748 14341 15804
rect 14341 15748 14397 15804
rect 14397 15748 14401 15804
rect 14337 15744 14401 15748
rect 14417 15804 14481 15808
rect 14417 15748 14421 15804
rect 14421 15748 14477 15804
rect 14477 15748 14481 15804
rect 14417 15744 14481 15748
rect 19467 15804 19531 15808
rect 19467 15748 19471 15804
rect 19471 15748 19527 15804
rect 19527 15748 19531 15804
rect 19467 15744 19531 15748
rect 19547 15804 19611 15808
rect 19547 15748 19551 15804
rect 19551 15748 19607 15804
rect 19607 15748 19611 15804
rect 19547 15744 19611 15748
rect 19627 15804 19691 15808
rect 19627 15748 19631 15804
rect 19631 15748 19687 15804
rect 19687 15748 19691 15804
rect 19627 15744 19691 15748
rect 19707 15804 19771 15808
rect 19707 15748 19711 15804
rect 19711 15748 19767 15804
rect 19767 15748 19771 15804
rect 19707 15744 19771 15748
rect 4257 15260 4321 15264
rect 4257 15204 4261 15260
rect 4261 15204 4317 15260
rect 4317 15204 4321 15260
rect 4257 15200 4321 15204
rect 4337 15260 4401 15264
rect 4337 15204 4341 15260
rect 4341 15204 4397 15260
rect 4397 15204 4401 15260
rect 4337 15200 4401 15204
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 9547 15260 9611 15264
rect 9547 15204 9551 15260
rect 9551 15204 9607 15260
rect 9607 15204 9611 15260
rect 9547 15200 9611 15204
rect 9627 15260 9691 15264
rect 9627 15204 9631 15260
rect 9631 15204 9687 15260
rect 9687 15204 9691 15260
rect 9627 15200 9691 15204
rect 9707 15260 9771 15264
rect 9707 15204 9711 15260
rect 9711 15204 9767 15260
rect 9767 15204 9771 15260
rect 9707 15200 9771 15204
rect 9787 15260 9851 15264
rect 9787 15204 9791 15260
rect 9791 15204 9847 15260
rect 9847 15204 9851 15260
rect 9787 15200 9851 15204
rect 14837 15260 14901 15264
rect 14837 15204 14841 15260
rect 14841 15204 14897 15260
rect 14897 15204 14901 15260
rect 14837 15200 14901 15204
rect 14917 15260 14981 15264
rect 14917 15204 14921 15260
rect 14921 15204 14977 15260
rect 14977 15204 14981 15260
rect 14917 15200 14981 15204
rect 14997 15260 15061 15264
rect 14997 15204 15001 15260
rect 15001 15204 15057 15260
rect 15057 15204 15061 15260
rect 14997 15200 15061 15204
rect 15077 15260 15141 15264
rect 15077 15204 15081 15260
rect 15081 15204 15137 15260
rect 15137 15204 15141 15260
rect 15077 15200 15141 15204
rect 20127 15260 20191 15264
rect 20127 15204 20131 15260
rect 20131 15204 20187 15260
rect 20187 15204 20191 15260
rect 20127 15200 20191 15204
rect 20207 15260 20271 15264
rect 20207 15204 20211 15260
rect 20211 15204 20267 15260
rect 20267 15204 20271 15260
rect 20207 15200 20271 15204
rect 20287 15260 20351 15264
rect 20287 15204 20291 15260
rect 20291 15204 20347 15260
rect 20347 15204 20351 15260
rect 20287 15200 20351 15204
rect 20367 15260 20431 15264
rect 20367 15204 20371 15260
rect 20371 15204 20427 15260
rect 20427 15204 20431 15260
rect 20367 15200 20431 15204
rect 3597 14716 3661 14720
rect 3597 14660 3601 14716
rect 3601 14660 3657 14716
rect 3657 14660 3661 14716
rect 3597 14656 3661 14660
rect 3677 14716 3741 14720
rect 3677 14660 3681 14716
rect 3681 14660 3737 14716
rect 3737 14660 3741 14716
rect 3677 14656 3741 14660
rect 3757 14716 3821 14720
rect 3757 14660 3761 14716
rect 3761 14660 3817 14716
rect 3817 14660 3821 14716
rect 3757 14656 3821 14660
rect 3837 14716 3901 14720
rect 3837 14660 3841 14716
rect 3841 14660 3897 14716
rect 3897 14660 3901 14716
rect 3837 14656 3901 14660
rect 8887 14716 8951 14720
rect 8887 14660 8891 14716
rect 8891 14660 8947 14716
rect 8947 14660 8951 14716
rect 8887 14656 8951 14660
rect 8967 14716 9031 14720
rect 8967 14660 8971 14716
rect 8971 14660 9027 14716
rect 9027 14660 9031 14716
rect 8967 14656 9031 14660
rect 9047 14716 9111 14720
rect 9047 14660 9051 14716
rect 9051 14660 9107 14716
rect 9107 14660 9111 14716
rect 9047 14656 9111 14660
rect 9127 14716 9191 14720
rect 9127 14660 9131 14716
rect 9131 14660 9187 14716
rect 9187 14660 9191 14716
rect 9127 14656 9191 14660
rect 14177 14716 14241 14720
rect 14177 14660 14181 14716
rect 14181 14660 14237 14716
rect 14237 14660 14241 14716
rect 14177 14656 14241 14660
rect 14257 14716 14321 14720
rect 14257 14660 14261 14716
rect 14261 14660 14317 14716
rect 14317 14660 14321 14716
rect 14257 14656 14321 14660
rect 14337 14716 14401 14720
rect 14337 14660 14341 14716
rect 14341 14660 14397 14716
rect 14397 14660 14401 14716
rect 14337 14656 14401 14660
rect 14417 14716 14481 14720
rect 14417 14660 14421 14716
rect 14421 14660 14477 14716
rect 14477 14660 14481 14716
rect 14417 14656 14481 14660
rect 19467 14716 19531 14720
rect 19467 14660 19471 14716
rect 19471 14660 19527 14716
rect 19527 14660 19531 14716
rect 19467 14656 19531 14660
rect 19547 14716 19611 14720
rect 19547 14660 19551 14716
rect 19551 14660 19607 14716
rect 19607 14660 19611 14716
rect 19547 14656 19611 14660
rect 19627 14716 19691 14720
rect 19627 14660 19631 14716
rect 19631 14660 19687 14716
rect 19687 14660 19691 14716
rect 19627 14656 19691 14660
rect 19707 14716 19771 14720
rect 19707 14660 19711 14716
rect 19711 14660 19767 14716
rect 19767 14660 19771 14716
rect 19707 14656 19771 14660
rect 4257 14172 4321 14176
rect 4257 14116 4261 14172
rect 4261 14116 4317 14172
rect 4317 14116 4321 14172
rect 4257 14112 4321 14116
rect 4337 14172 4401 14176
rect 4337 14116 4341 14172
rect 4341 14116 4397 14172
rect 4397 14116 4401 14172
rect 4337 14112 4401 14116
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 9547 14172 9611 14176
rect 9547 14116 9551 14172
rect 9551 14116 9607 14172
rect 9607 14116 9611 14172
rect 9547 14112 9611 14116
rect 9627 14172 9691 14176
rect 9627 14116 9631 14172
rect 9631 14116 9687 14172
rect 9687 14116 9691 14172
rect 9627 14112 9691 14116
rect 9707 14172 9771 14176
rect 9707 14116 9711 14172
rect 9711 14116 9767 14172
rect 9767 14116 9771 14172
rect 9707 14112 9771 14116
rect 9787 14172 9851 14176
rect 9787 14116 9791 14172
rect 9791 14116 9847 14172
rect 9847 14116 9851 14172
rect 9787 14112 9851 14116
rect 14837 14172 14901 14176
rect 14837 14116 14841 14172
rect 14841 14116 14897 14172
rect 14897 14116 14901 14172
rect 14837 14112 14901 14116
rect 14917 14172 14981 14176
rect 14917 14116 14921 14172
rect 14921 14116 14977 14172
rect 14977 14116 14981 14172
rect 14917 14112 14981 14116
rect 14997 14172 15061 14176
rect 14997 14116 15001 14172
rect 15001 14116 15057 14172
rect 15057 14116 15061 14172
rect 14997 14112 15061 14116
rect 15077 14172 15141 14176
rect 15077 14116 15081 14172
rect 15081 14116 15137 14172
rect 15137 14116 15141 14172
rect 15077 14112 15141 14116
rect 20127 14172 20191 14176
rect 20127 14116 20131 14172
rect 20131 14116 20187 14172
rect 20187 14116 20191 14172
rect 20127 14112 20191 14116
rect 20207 14172 20271 14176
rect 20207 14116 20211 14172
rect 20211 14116 20267 14172
rect 20267 14116 20271 14172
rect 20207 14112 20271 14116
rect 20287 14172 20351 14176
rect 20287 14116 20291 14172
rect 20291 14116 20347 14172
rect 20347 14116 20351 14172
rect 20287 14112 20351 14116
rect 20367 14172 20431 14176
rect 20367 14116 20371 14172
rect 20371 14116 20427 14172
rect 20427 14116 20431 14172
rect 20367 14112 20431 14116
rect 3597 13628 3661 13632
rect 3597 13572 3601 13628
rect 3601 13572 3657 13628
rect 3657 13572 3661 13628
rect 3597 13568 3661 13572
rect 3677 13628 3741 13632
rect 3677 13572 3681 13628
rect 3681 13572 3737 13628
rect 3737 13572 3741 13628
rect 3677 13568 3741 13572
rect 3757 13628 3821 13632
rect 3757 13572 3761 13628
rect 3761 13572 3817 13628
rect 3817 13572 3821 13628
rect 3757 13568 3821 13572
rect 3837 13628 3901 13632
rect 3837 13572 3841 13628
rect 3841 13572 3897 13628
rect 3897 13572 3901 13628
rect 3837 13568 3901 13572
rect 8887 13628 8951 13632
rect 8887 13572 8891 13628
rect 8891 13572 8947 13628
rect 8947 13572 8951 13628
rect 8887 13568 8951 13572
rect 8967 13628 9031 13632
rect 8967 13572 8971 13628
rect 8971 13572 9027 13628
rect 9027 13572 9031 13628
rect 8967 13568 9031 13572
rect 9047 13628 9111 13632
rect 9047 13572 9051 13628
rect 9051 13572 9107 13628
rect 9107 13572 9111 13628
rect 9047 13568 9111 13572
rect 9127 13628 9191 13632
rect 9127 13572 9131 13628
rect 9131 13572 9187 13628
rect 9187 13572 9191 13628
rect 9127 13568 9191 13572
rect 14177 13628 14241 13632
rect 14177 13572 14181 13628
rect 14181 13572 14237 13628
rect 14237 13572 14241 13628
rect 14177 13568 14241 13572
rect 14257 13628 14321 13632
rect 14257 13572 14261 13628
rect 14261 13572 14317 13628
rect 14317 13572 14321 13628
rect 14257 13568 14321 13572
rect 14337 13628 14401 13632
rect 14337 13572 14341 13628
rect 14341 13572 14397 13628
rect 14397 13572 14401 13628
rect 14337 13568 14401 13572
rect 14417 13628 14481 13632
rect 14417 13572 14421 13628
rect 14421 13572 14477 13628
rect 14477 13572 14481 13628
rect 14417 13568 14481 13572
rect 19467 13628 19531 13632
rect 19467 13572 19471 13628
rect 19471 13572 19527 13628
rect 19527 13572 19531 13628
rect 19467 13568 19531 13572
rect 19547 13628 19611 13632
rect 19547 13572 19551 13628
rect 19551 13572 19607 13628
rect 19607 13572 19611 13628
rect 19547 13568 19611 13572
rect 19627 13628 19691 13632
rect 19627 13572 19631 13628
rect 19631 13572 19687 13628
rect 19687 13572 19691 13628
rect 19627 13568 19691 13572
rect 19707 13628 19771 13632
rect 19707 13572 19711 13628
rect 19711 13572 19767 13628
rect 19767 13572 19771 13628
rect 19707 13568 19771 13572
rect 4257 13084 4321 13088
rect 4257 13028 4261 13084
rect 4261 13028 4317 13084
rect 4317 13028 4321 13084
rect 4257 13024 4321 13028
rect 4337 13084 4401 13088
rect 4337 13028 4341 13084
rect 4341 13028 4397 13084
rect 4397 13028 4401 13084
rect 4337 13024 4401 13028
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 9547 13084 9611 13088
rect 9547 13028 9551 13084
rect 9551 13028 9607 13084
rect 9607 13028 9611 13084
rect 9547 13024 9611 13028
rect 9627 13084 9691 13088
rect 9627 13028 9631 13084
rect 9631 13028 9687 13084
rect 9687 13028 9691 13084
rect 9627 13024 9691 13028
rect 9707 13084 9771 13088
rect 9707 13028 9711 13084
rect 9711 13028 9767 13084
rect 9767 13028 9771 13084
rect 9707 13024 9771 13028
rect 9787 13084 9851 13088
rect 9787 13028 9791 13084
rect 9791 13028 9847 13084
rect 9847 13028 9851 13084
rect 9787 13024 9851 13028
rect 14837 13084 14901 13088
rect 14837 13028 14841 13084
rect 14841 13028 14897 13084
rect 14897 13028 14901 13084
rect 14837 13024 14901 13028
rect 14917 13084 14981 13088
rect 14917 13028 14921 13084
rect 14921 13028 14977 13084
rect 14977 13028 14981 13084
rect 14917 13024 14981 13028
rect 14997 13084 15061 13088
rect 14997 13028 15001 13084
rect 15001 13028 15057 13084
rect 15057 13028 15061 13084
rect 14997 13024 15061 13028
rect 15077 13084 15141 13088
rect 15077 13028 15081 13084
rect 15081 13028 15137 13084
rect 15137 13028 15141 13084
rect 15077 13024 15141 13028
rect 20127 13084 20191 13088
rect 20127 13028 20131 13084
rect 20131 13028 20187 13084
rect 20187 13028 20191 13084
rect 20127 13024 20191 13028
rect 20207 13084 20271 13088
rect 20207 13028 20211 13084
rect 20211 13028 20267 13084
rect 20267 13028 20271 13084
rect 20207 13024 20271 13028
rect 20287 13084 20351 13088
rect 20287 13028 20291 13084
rect 20291 13028 20347 13084
rect 20347 13028 20351 13084
rect 20287 13024 20351 13028
rect 20367 13084 20431 13088
rect 20367 13028 20371 13084
rect 20371 13028 20427 13084
rect 20427 13028 20431 13084
rect 20367 13024 20431 13028
rect 3597 12540 3661 12544
rect 3597 12484 3601 12540
rect 3601 12484 3657 12540
rect 3657 12484 3661 12540
rect 3597 12480 3661 12484
rect 3677 12540 3741 12544
rect 3677 12484 3681 12540
rect 3681 12484 3737 12540
rect 3737 12484 3741 12540
rect 3677 12480 3741 12484
rect 3757 12540 3821 12544
rect 3757 12484 3761 12540
rect 3761 12484 3817 12540
rect 3817 12484 3821 12540
rect 3757 12480 3821 12484
rect 3837 12540 3901 12544
rect 3837 12484 3841 12540
rect 3841 12484 3897 12540
rect 3897 12484 3901 12540
rect 3837 12480 3901 12484
rect 8887 12540 8951 12544
rect 8887 12484 8891 12540
rect 8891 12484 8947 12540
rect 8947 12484 8951 12540
rect 8887 12480 8951 12484
rect 8967 12540 9031 12544
rect 8967 12484 8971 12540
rect 8971 12484 9027 12540
rect 9027 12484 9031 12540
rect 8967 12480 9031 12484
rect 9047 12540 9111 12544
rect 9047 12484 9051 12540
rect 9051 12484 9107 12540
rect 9107 12484 9111 12540
rect 9047 12480 9111 12484
rect 9127 12540 9191 12544
rect 9127 12484 9131 12540
rect 9131 12484 9187 12540
rect 9187 12484 9191 12540
rect 9127 12480 9191 12484
rect 14177 12540 14241 12544
rect 14177 12484 14181 12540
rect 14181 12484 14237 12540
rect 14237 12484 14241 12540
rect 14177 12480 14241 12484
rect 14257 12540 14321 12544
rect 14257 12484 14261 12540
rect 14261 12484 14317 12540
rect 14317 12484 14321 12540
rect 14257 12480 14321 12484
rect 14337 12540 14401 12544
rect 14337 12484 14341 12540
rect 14341 12484 14397 12540
rect 14397 12484 14401 12540
rect 14337 12480 14401 12484
rect 14417 12540 14481 12544
rect 14417 12484 14421 12540
rect 14421 12484 14477 12540
rect 14477 12484 14481 12540
rect 14417 12480 14481 12484
rect 19467 12540 19531 12544
rect 19467 12484 19471 12540
rect 19471 12484 19527 12540
rect 19527 12484 19531 12540
rect 19467 12480 19531 12484
rect 19547 12540 19611 12544
rect 19547 12484 19551 12540
rect 19551 12484 19607 12540
rect 19607 12484 19611 12540
rect 19547 12480 19611 12484
rect 19627 12540 19691 12544
rect 19627 12484 19631 12540
rect 19631 12484 19687 12540
rect 19687 12484 19691 12540
rect 19627 12480 19691 12484
rect 19707 12540 19771 12544
rect 19707 12484 19711 12540
rect 19711 12484 19767 12540
rect 19767 12484 19771 12540
rect 19707 12480 19771 12484
rect 4257 11996 4321 12000
rect 4257 11940 4261 11996
rect 4261 11940 4317 11996
rect 4317 11940 4321 11996
rect 4257 11936 4321 11940
rect 4337 11996 4401 12000
rect 4337 11940 4341 11996
rect 4341 11940 4397 11996
rect 4397 11940 4401 11996
rect 4337 11936 4401 11940
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 9547 11996 9611 12000
rect 9547 11940 9551 11996
rect 9551 11940 9607 11996
rect 9607 11940 9611 11996
rect 9547 11936 9611 11940
rect 9627 11996 9691 12000
rect 9627 11940 9631 11996
rect 9631 11940 9687 11996
rect 9687 11940 9691 11996
rect 9627 11936 9691 11940
rect 9707 11996 9771 12000
rect 9707 11940 9711 11996
rect 9711 11940 9767 11996
rect 9767 11940 9771 11996
rect 9707 11936 9771 11940
rect 9787 11996 9851 12000
rect 9787 11940 9791 11996
rect 9791 11940 9847 11996
rect 9847 11940 9851 11996
rect 9787 11936 9851 11940
rect 14837 11996 14901 12000
rect 14837 11940 14841 11996
rect 14841 11940 14897 11996
rect 14897 11940 14901 11996
rect 14837 11936 14901 11940
rect 14917 11996 14981 12000
rect 14917 11940 14921 11996
rect 14921 11940 14977 11996
rect 14977 11940 14981 11996
rect 14917 11936 14981 11940
rect 14997 11996 15061 12000
rect 14997 11940 15001 11996
rect 15001 11940 15057 11996
rect 15057 11940 15061 11996
rect 14997 11936 15061 11940
rect 15077 11996 15141 12000
rect 15077 11940 15081 11996
rect 15081 11940 15137 11996
rect 15137 11940 15141 11996
rect 15077 11936 15141 11940
rect 20127 11996 20191 12000
rect 20127 11940 20131 11996
rect 20131 11940 20187 11996
rect 20187 11940 20191 11996
rect 20127 11936 20191 11940
rect 20207 11996 20271 12000
rect 20207 11940 20211 11996
rect 20211 11940 20267 11996
rect 20267 11940 20271 11996
rect 20207 11936 20271 11940
rect 20287 11996 20351 12000
rect 20287 11940 20291 11996
rect 20291 11940 20347 11996
rect 20347 11940 20351 11996
rect 20287 11936 20351 11940
rect 20367 11996 20431 12000
rect 20367 11940 20371 11996
rect 20371 11940 20427 11996
rect 20427 11940 20431 11996
rect 20367 11936 20431 11940
rect 3597 11452 3661 11456
rect 3597 11396 3601 11452
rect 3601 11396 3657 11452
rect 3657 11396 3661 11452
rect 3597 11392 3661 11396
rect 3677 11452 3741 11456
rect 3677 11396 3681 11452
rect 3681 11396 3737 11452
rect 3737 11396 3741 11452
rect 3677 11392 3741 11396
rect 3757 11452 3821 11456
rect 3757 11396 3761 11452
rect 3761 11396 3817 11452
rect 3817 11396 3821 11452
rect 3757 11392 3821 11396
rect 3837 11452 3901 11456
rect 3837 11396 3841 11452
rect 3841 11396 3897 11452
rect 3897 11396 3901 11452
rect 3837 11392 3901 11396
rect 8887 11452 8951 11456
rect 8887 11396 8891 11452
rect 8891 11396 8947 11452
rect 8947 11396 8951 11452
rect 8887 11392 8951 11396
rect 8967 11452 9031 11456
rect 8967 11396 8971 11452
rect 8971 11396 9027 11452
rect 9027 11396 9031 11452
rect 8967 11392 9031 11396
rect 9047 11452 9111 11456
rect 9047 11396 9051 11452
rect 9051 11396 9107 11452
rect 9107 11396 9111 11452
rect 9047 11392 9111 11396
rect 9127 11452 9191 11456
rect 9127 11396 9131 11452
rect 9131 11396 9187 11452
rect 9187 11396 9191 11452
rect 9127 11392 9191 11396
rect 14177 11452 14241 11456
rect 14177 11396 14181 11452
rect 14181 11396 14237 11452
rect 14237 11396 14241 11452
rect 14177 11392 14241 11396
rect 14257 11452 14321 11456
rect 14257 11396 14261 11452
rect 14261 11396 14317 11452
rect 14317 11396 14321 11452
rect 14257 11392 14321 11396
rect 14337 11452 14401 11456
rect 14337 11396 14341 11452
rect 14341 11396 14397 11452
rect 14397 11396 14401 11452
rect 14337 11392 14401 11396
rect 14417 11452 14481 11456
rect 14417 11396 14421 11452
rect 14421 11396 14477 11452
rect 14477 11396 14481 11452
rect 14417 11392 14481 11396
rect 19467 11452 19531 11456
rect 19467 11396 19471 11452
rect 19471 11396 19527 11452
rect 19527 11396 19531 11452
rect 19467 11392 19531 11396
rect 19547 11452 19611 11456
rect 19547 11396 19551 11452
rect 19551 11396 19607 11452
rect 19607 11396 19611 11452
rect 19547 11392 19611 11396
rect 19627 11452 19691 11456
rect 19627 11396 19631 11452
rect 19631 11396 19687 11452
rect 19687 11396 19691 11452
rect 19627 11392 19691 11396
rect 19707 11452 19771 11456
rect 19707 11396 19711 11452
rect 19711 11396 19767 11452
rect 19767 11396 19771 11452
rect 19707 11392 19771 11396
rect 4257 10908 4321 10912
rect 4257 10852 4261 10908
rect 4261 10852 4317 10908
rect 4317 10852 4321 10908
rect 4257 10848 4321 10852
rect 4337 10908 4401 10912
rect 4337 10852 4341 10908
rect 4341 10852 4397 10908
rect 4397 10852 4401 10908
rect 4337 10848 4401 10852
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 9547 10908 9611 10912
rect 9547 10852 9551 10908
rect 9551 10852 9607 10908
rect 9607 10852 9611 10908
rect 9547 10848 9611 10852
rect 9627 10908 9691 10912
rect 9627 10852 9631 10908
rect 9631 10852 9687 10908
rect 9687 10852 9691 10908
rect 9627 10848 9691 10852
rect 9707 10908 9771 10912
rect 9707 10852 9711 10908
rect 9711 10852 9767 10908
rect 9767 10852 9771 10908
rect 9707 10848 9771 10852
rect 9787 10908 9851 10912
rect 9787 10852 9791 10908
rect 9791 10852 9847 10908
rect 9847 10852 9851 10908
rect 9787 10848 9851 10852
rect 14837 10908 14901 10912
rect 14837 10852 14841 10908
rect 14841 10852 14897 10908
rect 14897 10852 14901 10908
rect 14837 10848 14901 10852
rect 14917 10908 14981 10912
rect 14917 10852 14921 10908
rect 14921 10852 14977 10908
rect 14977 10852 14981 10908
rect 14917 10848 14981 10852
rect 14997 10908 15061 10912
rect 14997 10852 15001 10908
rect 15001 10852 15057 10908
rect 15057 10852 15061 10908
rect 14997 10848 15061 10852
rect 15077 10908 15141 10912
rect 15077 10852 15081 10908
rect 15081 10852 15137 10908
rect 15137 10852 15141 10908
rect 15077 10848 15141 10852
rect 20127 10908 20191 10912
rect 20127 10852 20131 10908
rect 20131 10852 20187 10908
rect 20187 10852 20191 10908
rect 20127 10848 20191 10852
rect 20207 10908 20271 10912
rect 20207 10852 20211 10908
rect 20211 10852 20267 10908
rect 20267 10852 20271 10908
rect 20207 10848 20271 10852
rect 20287 10908 20351 10912
rect 20287 10852 20291 10908
rect 20291 10852 20347 10908
rect 20347 10852 20351 10908
rect 20287 10848 20351 10852
rect 20367 10908 20431 10912
rect 20367 10852 20371 10908
rect 20371 10852 20427 10908
rect 20427 10852 20431 10908
rect 20367 10848 20431 10852
rect 3597 10364 3661 10368
rect 3597 10308 3601 10364
rect 3601 10308 3657 10364
rect 3657 10308 3661 10364
rect 3597 10304 3661 10308
rect 3677 10364 3741 10368
rect 3677 10308 3681 10364
rect 3681 10308 3737 10364
rect 3737 10308 3741 10364
rect 3677 10304 3741 10308
rect 3757 10364 3821 10368
rect 3757 10308 3761 10364
rect 3761 10308 3817 10364
rect 3817 10308 3821 10364
rect 3757 10304 3821 10308
rect 3837 10364 3901 10368
rect 3837 10308 3841 10364
rect 3841 10308 3897 10364
rect 3897 10308 3901 10364
rect 3837 10304 3901 10308
rect 8887 10364 8951 10368
rect 8887 10308 8891 10364
rect 8891 10308 8947 10364
rect 8947 10308 8951 10364
rect 8887 10304 8951 10308
rect 8967 10364 9031 10368
rect 8967 10308 8971 10364
rect 8971 10308 9027 10364
rect 9027 10308 9031 10364
rect 8967 10304 9031 10308
rect 9047 10364 9111 10368
rect 9047 10308 9051 10364
rect 9051 10308 9107 10364
rect 9107 10308 9111 10364
rect 9047 10304 9111 10308
rect 9127 10364 9191 10368
rect 9127 10308 9131 10364
rect 9131 10308 9187 10364
rect 9187 10308 9191 10364
rect 9127 10304 9191 10308
rect 14177 10364 14241 10368
rect 14177 10308 14181 10364
rect 14181 10308 14237 10364
rect 14237 10308 14241 10364
rect 14177 10304 14241 10308
rect 14257 10364 14321 10368
rect 14257 10308 14261 10364
rect 14261 10308 14317 10364
rect 14317 10308 14321 10364
rect 14257 10304 14321 10308
rect 14337 10364 14401 10368
rect 14337 10308 14341 10364
rect 14341 10308 14397 10364
rect 14397 10308 14401 10364
rect 14337 10304 14401 10308
rect 14417 10364 14481 10368
rect 14417 10308 14421 10364
rect 14421 10308 14477 10364
rect 14477 10308 14481 10364
rect 14417 10304 14481 10308
rect 19467 10364 19531 10368
rect 19467 10308 19471 10364
rect 19471 10308 19527 10364
rect 19527 10308 19531 10364
rect 19467 10304 19531 10308
rect 19547 10364 19611 10368
rect 19547 10308 19551 10364
rect 19551 10308 19607 10364
rect 19607 10308 19611 10364
rect 19547 10304 19611 10308
rect 19627 10364 19691 10368
rect 19627 10308 19631 10364
rect 19631 10308 19687 10364
rect 19687 10308 19691 10364
rect 19627 10304 19691 10308
rect 19707 10364 19771 10368
rect 19707 10308 19711 10364
rect 19711 10308 19767 10364
rect 19767 10308 19771 10364
rect 19707 10304 19771 10308
rect 4257 9820 4321 9824
rect 4257 9764 4261 9820
rect 4261 9764 4317 9820
rect 4317 9764 4321 9820
rect 4257 9760 4321 9764
rect 4337 9820 4401 9824
rect 4337 9764 4341 9820
rect 4341 9764 4397 9820
rect 4397 9764 4401 9820
rect 4337 9760 4401 9764
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 9547 9820 9611 9824
rect 9547 9764 9551 9820
rect 9551 9764 9607 9820
rect 9607 9764 9611 9820
rect 9547 9760 9611 9764
rect 9627 9820 9691 9824
rect 9627 9764 9631 9820
rect 9631 9764 9687 9820
rect 9687 9764 9691 9820
rect 9627 9760 9691 9764
rect 9707 9820 9771 9824
rect 9707 9764 9711 9820
rect 9711 9764 9767 9820
rect 9767 9764 9771 9820
rect 9707 9760 9771 9764
rect 9787 9820 9851 9824
rect 9787 9764 9791 9820
rect 9791 9764 9847 9820
rect 9847 9764 9851 9820
rect 9787 9760 9851 9764
rect 14837 9820 14901 9824
rect 14837 9764 14841 9820
rect 14841 9764 14897 9820
rect 14897 9764 14901 9820
rect 14837 9760 14901 9764
rect 14917 9820 14981 9824
rect 14917 9764 14921 9820
rect 14921 9764 14977 9820
rect 14977 9764 14981 9820
rect 14917 9760 14981 9764
rect 14997 9820 15061 9824
rect 14997 9764 15001 9820
rect 15001 9764 15057 9820
rect 15057 9764 15061 9820
rect 14997 9760 15061 9764
rect 15077 9820 15141 9824
rect 15077 9764 15081 9820
rect 15081 9764 15137 9820
rect 15137 9764 15141 9820
rect 15077 9760 15141 9764
rect 20127 9820 20191 9824
rect 20127 9764 20131 9820
rect 20131 9764 20187 9820
rect 20187 9764 20191 9820
rect 20127 9760 20191 9764
rect 20207 9820 20271 9824
rect 20207 9764 20211 9820
rect 20211 9764 20267 9820
rect 20267 9764 20271 9820
rect 20207 9760 20271 9764
rect 20287 9820 20351 9824
rect 20287 9764 20291 9820
rect 20291 9764 20347 9820
rect 20347 9764 20351 9820
rect 20287 9760 20351 9764
rect 20367 9820 20431 9824
rect 20367 9764 20371 9820
rect 20371 9764 20427 9820
rect 20427 9764 20431 9820
rect 20367 9760 20431 9764
rect 3597 9276 3661 9280
rect 3597 9220 3601 9276
rect 3601 9220 3657 9276
rect 3657 9220 3661 9276
rect 3597 9216 3661 9220
rect 3677 9276 3741 9280
rect 3677 9220 3681 9276
rect 3681 9220 3737 9276
rect 3737 9220 3741 9276
rect 3677 9216 3741 9220
rect 3757 9276 3821 9280
rect 3757 9220 3761 9276
rect 3761 9220 3817 9276
rect 3817 9220 3821 9276
rect 3757 9216 3821 9220
rect 3837 9276 3901 9280
rect 3837 9220 3841 9276
rect 3841 9220 3897 9276
rect 3897 9220 3901 9276
rect 3837 9216 3901 9220
rect 8887 9276 8951 9280
rect 8887 9220 8891 9276
rect 8891 9220 8947 9276
rect 8947 9220 8951 9276
rect 8887 9216 8951 9220
rect 8967 9276 9031 9280
rect 8967 9220 8971 9276
rect 8971 9220 9027 9276
rect 9027 9220 9031 9276
rect 8967 9216 9031 9220
rect 9047 9276 9111 9280
rect 9047 9220 9051 9276
rect 9051 9220 9107 9276
rect 9107 9220 9111 9276
rect 9047 9216 9111 9220
rect 9127 9276 9191 9280
rect 9127 9220 9131 9276
rect 9131 9220 9187 9276
rect 9187 9220 9191 9276
rect 9127 9216 9191 9220
rect 14177 9276 14241 9280
rect 14177 9220 14181 9276
rect 14181 9220 14237 9276
rect 14237 9220 14241 9276
rect 14177 9216 14241 9220
rect 14257 9276 14321 9280
rect 14257 9220 14261 9276
rect 14261 9220 14317 9276
rect 14317 9220 14321 9276
rect 14257 9216 14321 9220
rect 14337 9276 14401 9280
rect 14337 9220 14341 9276
rect 14341 9220 14397 9276
rect 14397 9220 14401 9276
rect 14337 9216 14401 9220
rect 14417 9276 14481 9280
rect 14417 9220 14421 9276
rect 14421 9220 14477 9276
rect 14477 9220 14481 9276
rect 14417 9216 14481 9220
rect 19467 9276 19531 9280
rect 19467 9220 19471 9276
rect 19471 9220 19527 9276
rect 19527 9220 19531 9276
rect 19467 9216 19531 9220
rect 19547 9276 19611 9280
rect 19547 9220 19551 9276
rect 19551 9220 19607 9276
rect 19607 9220 19611 9276
rect 19547 9216 19611 9220
rect 19627 9276 19691 9280
rect 19627 9220 19631 9276
rect 19631 9220 19687 9276
rect 19687 9220 19691 9276
rect 19627 9216 19691 9220
rect 19707 9276 19771 9280
rect 19707 9220 19711 9276
rect 19711 9220 19767 9276
rect 19767 9220 19771 9276
rect 19707 9216 19771 9220
rect 4257 8732 4321 8736
rect 4257 8676 4261 8732
rect 4261 8676 4317 8732
rect 4317 8676 4321 8732
rect 4257 8672 4321 8676
rect 4337 8732 4401 8736
rect 4337 8676 4341 8732
rect 4341 8676 4397 8732
rect 4397 8676 4401 8732
rect 4337 8672 4401 8676
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 9547 8732 9611 8736
rect 9547 8676 9551 8732
rect 9551 8676 9607 8732
rect 9607 8676 9611 8732
rect 9547 8672 9611 8676
rect 9627 8732 9691 8736
rect 9627 8676 9631 8732
rect 9631 8676 9687 8732
rect 9687 8676 9691 8732
rect 9627 8672 9691 8676
rect 9707 8732 9771 8736
rect 9707 8676 9711 8732
rect 9711 8676 9767 8732
rect 9767 8676 9771 8732
rect 9707 8672 9771 8676
rect 9787 8732 9851 8736
rect 9787 8676 9791 8732
rect 9791 8676 9847 8732
rect 9847 8676 9851 8732
rect 9787 8672 9851 8676
rect 14837 8732 14901 8736
rect 14837 8676 14841 8732
rect 14841 8676 14897 8732
rect 14897 8676 14901 8732
rect 14837 8672 14901 8676
rect 14917 8732 14981 8736
rect 14917 8676 14921 8732
rect 14921 8676 14977 8732
rect 14977 8676 14981 8732
rect 14917 8672 14981 8676
rect 14997 8732 15061 8736
rect 14997 8676 15001 8732
rect 15001 8676 15057 8732
rect 15057 8676 15061 8732
rect 14997 8672 15061 8676
rect 15077 8732 15141 8736
rect 15077 8676 15081 8732
rect 15081 8676 15137 8732
rect 15137 8676 15141 8732
rect 15077 8672 15141 8676
rect 20127 8732 20191 8736
rect 20127 8676 20131 8732
rect 20131 8676 20187 8732
rect 20187 8676 20191 8732
rect 20127 8672 20191 8676
rect 20207 8732 20271 8736
rect 20207 8676 20211 8732
rect 20211 8676 20267 8732
rect 20267 8676 20271 8732
rect 20207 8672 20271 8676
rect 20287 8732 20351 8736
rect 20287 8676 20291 8732
rect 20291 8676 20347 8732
rect 20347 8676 20351 8732
rect 20287 8672 20351 8676
rect 20367 8732 20431 8736
rect 20367 8676 20371 8732
rect 20371 8676 20427 8732
rect 20427 8676 20431 8732
rect 20367 8672 20431 8676
rect 3597 8188 3661 8192
rect 3597 8132 3601 8188
rect 3601 8132 3657 8188
rect 3657 8132 3661 8188
rect 3597 8128 3661 8132
rect 3677 8188 3741 8192
rect 3677 8132 3681 8188
rect 3681 8132 3737 8188
rect 3737 8132 3741 8188
rect 3677 8128 3741 8132
rect 3757 8188 3821 8192
rect 3757 8132 3761 8188
rect 3761 8132 3817 8188
rect 3817 8132 3821 8188
rect 3757 8128 3821 8132
rect 3837 8188 3901 8192
rect 3837 8132 3841 8188
rect 3841 8132 3897 8188
rect 3897 8132 3901 8188
rect 3837 8128 3901 8132
rect 8887 8188 8951 8192
rect 8887 8132 8891 8188
rect 8891 8132 8947 8188
rect 8947 8132 8951 8188
rect 8887 8128 8951 8132
rect 8967 8188 9031 8192
rect 8967 8132 8971 8188
rect 8971 8132 9027 8188
rect 9027 8132 9031 8188
rect 8967 8128 9031 8132
rect 9047 8188 9111 8192
rect 9047 8132 9051 8188
rect 9051 8132 9107 8188
rect 9107 8132 9111 8188
rect 9047 8128 9111 8132
rect 9127 8188 9191 8192
rect 9127 8132 9131 8188
rect 9131 8132 9187 8188
rect 9187 8132 9191 8188
rect 9127 8128 9191 8132
rect 14177 8188 14241 8192
rect 14177 8132 14181 8188
rect 14181 8132 14237 8188
rect 14237 8132 14241 8188
rect 14177 8128 14241 8132
rect 14257 8188 14321 8192
rect 14257 8132 14261 8188
rect 14261 8132 14317 8188
rect 14317 8132 14321 8188
rect 14257 8128 14321 8132
rect 14337 8188 14401 8192
rect 14337 8132 14341 8188
rect 14341 8132 14397 8188
rect 14397 8132 14401 8188
rect 14337 8128 14401 8132
rect 14417 8188 14481 8192
rect 14417 8132 14421 8188
rect 14421 8132 14477 8188
rect 14477 8132 14481 8188
rect 14417 8128 14481 8132
rect 19467 8188 19531 8192
rect 19467 8132 19471 8188
rect 19471 8132 19527 8188
rect 19527 8132 19531 8188
rect 19467 8128 19531 8132
rect 19547 8188 19611 8192
rect 19547 8132 19551 8188
rect 19551 8132 19607 8188
rect 19607 8132 19611 8188
rect 19547 8128 19611 8132
rect 19627 8188 19691 8192
rect 19627 8132 19631 8188
rect 19631 8132 19687 8188
rect 19687 8132 19691 8188
rect 19627 8128 19691 8132
rect 19707 8188 19771 8192
rect 19707 8132 19711 8188
rect 19711 8132 19767 8188
rect 19767 8132 19771 8188
rect 19707 8128 19771 8132
rect 4257 7644 4321 7648
rect 4257 7588 4261 7644
rect 4261 7588 4317 7644
rect 4317 7588 4321 7644
rect 4257 7584 4321 7588
rect 4337 7644 4401 7648
rect 4337 7588 4341 7644
rect 4341 7588 4397 7644
rect 4397 7588 4401 7644
rect 4337 7584 4401 7588
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 9547 7644 9611 7648
rect 9547 7588 9551 7644
rect 9551 7588 9607 7644
rect 9607 7588 9611 7644
rect 9547 7584 9611 7588
rect 9627 7644 9691 7648
rect 9627 7588 9631 7644
rect 9631 7588 9687 7644
rect 9687 7588 9691 7644
rect 9627 7584 9691 7588
rect 9707 7644 9771 7648
rect 9707 7588 9711 7644
rect 9711 7588 9767 7644
rect 9767 7588 9771 7644
rect 9707 7584 9771 7588
rect 9787 7644 9851 7648
rect 9787 7588 9791 7644
rect 9791 7588 9847 7644
rect 9847 7588 9851 7644
rect 9787 7584 9851 7588
rect 14837 7644 14901 7648
rect 14837 7588 14841 7644
rect 14841 7588 14897 7644
rect 14897 7588 14901 7644
rect 14837 7584 14901 7588
rect 14917 7644 14981 7648
rect 14917 7588 14921 7644
rect 14921 7588 14977 7644
rect 14977 7588 14981 7644
rect 14917 7584 14981 7588
rect 14997 7644 15061 7648
rect 14997 7588 15001 7644
rect 15001 7588 15057 7644
rect 15057 7588 15061 7644
rect 14997 7584 15061 7588
rect 15077 7644 15141 7648
rect 15077 7588 15081 7644
rect 15081 7588 15137 7644
rect 15137 7588 15141 7644
rect 15077 7584 15141 7588
rect 20127 7644 20191 7648
rect 20127 7588 20131 7644
rect 20131 7588 20187 7644
rect 20187 7588 20191 7644
rect 20127 7584 20191 7588
rect 20207 7644 20271 7648
rect 20207 7588 20211 7644
rect 20211 7588 20267 7644
rect 20267 7588 20271 7644
rect 20207 7584 20271 7588
rect 20287 7644 20351 7648
rect 20287 7588 20291 7644
rect 20291 7588 20347 7644
rect 20347 7588 20351 7644
rect 20287 7584 20351 7588
rect 20367 7644 20431 7648
rect 20367 7588 20371 7644
rect 20371 7588 20427 7644
rect 20427 7588 20431 7644
rect 20367 7584 20431 7588
rect 3597 7100 3661 7104
rect 3597 7044 3601 7100
rect 3601 7044 3657 7100
rect 3657 7044 3661 7100
rect 3597 7040 3661 7044
rect 3677 7100 3741 7104
rect 3677 7044 3681 7100
rect 3681 7044 3737 7100
rect 3737 7044 3741 7100
rect 3677 7040 3741 7044
rect 3757 7100 3821 7104
rect 3757 7044 3761 7100
rect 3761 7044 3817 7100
rect 3817 7044 3821 7100
rect 3757 7040 3821 7044
rect 3837 7100 3901 7104
rect 3837 7044 3841 7100
rect 3841 7044 3897 7100
rect 3897 7044 3901 7100
rect 3837 7040 3901 7044
rect 8887 7100 8951 7104
rect 8887 7044 8891 7100
rect 8891 7044 8947 7100
rect 8947 7044 8951 7100
rect 8887 7040 8951 7044
rect 8967 7100 9031 7104
rect 8967 7044 8971 7100
rect 8971 7044 9027 7100
rect 9027 7044 9031 7100
rect 8967 7040 9031 7044
rect 9047 7100 9111 7104
rect 9047 7044 9051 7100
rect 9051 7044 9107 7100
rect 9107 7044 9111 7100
rect 9047 7040 9111 7044
rect 9127 7100 9191 7104
rect 9127 7044 9131 7100
rect 9131 7044 9187 7100
rect 9187 7044 9191 7100
rect 9127 7040 9191 7044
rect 14177 7100 14241 7104
rect 14177 7044 14181 7100
rect 14181 7044 14237 7100
rect 14237 7044 14241 7100
rect 14177 7040 14241 7044
rect 14257 7100 14321 7104
rect 14257 7044 14261 7100
rect 14261 7044 14317 7100
rect 14317 7044 14321 7100
rect 14257 7040 14321 7044
rect 14337 7100 14401 7104
rect 14337 7044 14341 7100
rect 14341 7044 14397 7100
rect 14397 7044 14401 7100
rect 14337 7040 14401 7044
rect 14417 7100 14481 7104
rect 14417 7044 14421 7100
rect 14421 7044 14477 7100
rect 14477 7044 14481 7100
rect 14417 7040 14481 7044
rect 19467 7100 19531 7104
rect 19467 7044 19471 7100
rect 19471 7044 19527 7100
rect 19527 7044 19531 7100
rect 19467 7040 19531 7044
rect 19547 7100 19611 7104
rect 19547 7044 19551 7100
rect 19551 7044 19607 7100
rect 19607 7044 19611 7100
rect 19547 7040 19611 7044
rect 19627 7100 19691 7104
rect 19627 7044 19631 7100
rect 19631 7044 19687 7100
rect 19687 7044 19691 7100
rect 19627 7040 19691 7044
rect 19707 7100 19771 7104
rect 19707 7044 19711 7100
rect 19711 7044 19767 7100
rect 19767 7044 19771 7100
rect 19707 7040 19771 7044
rect 4257 6556 4321 6560
rect 4257 6500 4261 6556
rect 4261 6500 4317 6556
rect 4317 6500 4321 6556
rect 4257 6496 4321 6500
rect 4337 6556 4401 6560
rect 4337 6500 4341 6556
rect 4341 6500 4397 6556
rect 4397 6500 4401 6556
rect 4337 6496 4401 6500
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 9547 6556 9611 6560
rect 9547 6500 9551 6556
rect 9551 6500 9607 6556
rect 9607 6500 9611 6556
rect 9547 6496 9611 6500
rect 9627 6556 9691 6560
rect 9627 6500 9631 6556
rect 9631 6500 9687 6556
rect 9687 6500 9691 6556
rect 9627 6496 9691 6500
rect 9707 6556 9771 6560
rect 9707 6500 9711 6556
rect 9711 6500 9767 6556
rect 9767 6500 9771 6556
rect 9707 6496 9771 6500
rect 9787 6556 9851 6560
rect 9787 6500 9791 6556
rect 9791 6500 9847 6556
rect 9847 6500 9851 6556
rect 9787 6496 9851 6500
rect 14837 6556 14901 6560
rect 14837 6500 14841 6556
rect 14841 6500 14897 6556
rect 14897 6500 14901 6556
rect 14837 6496 14901 6500
rect 14917 6556 14981 6560
rect 14917 6500 14921 6556
rect 14921 6500 14977 6556
rect 14977 6500 14981 6556
rect 14917 6496 14981 6500
rect 14997 6556 15061 6560
rect 14997 6500 15001 6556
rect 15001 6500 15057 6556
rect 15057 6500 15061 6556
rect 14997 6496 15061 6500
rect 15077 6556 15141 6560
rect 15077 6500 15081 6556
rect 15081 6500 15137 6556
rect 15137 6500 15141 6556
rect 15077 6496 15141 6500
rect 20127 6556 20191 6560
rect 20127 6500 20131 6556
rect 20131 6500 20187 6556
rect 20187 6500 20191 6556
rect 20127 6496 20191 6500
rect 20207 6556 20271 6560
rect 20207 6500 20211 6556
rect 20211 6500 20267 6556
rect 20267 6500 20271 6556
rect 20207 6496 20271 6500
rect 20287 6556 20351 6560
rect 20287 6500 20291 6556
rect 20291 6500 20347 6556
rect 20347 6500 20351 6556
rect 20287 6496 20351 6500
rect 20367 6556 20431 6560
rect 20367 6500 20371 6556
rect 20371 6500 20427 6556
rect 20427 6500 20431 6556
rect 20367 6496 20431 6500
rect 3597 6012 3661 6016
rect 3597 5956 3601 6012
rect 3601 5956 3657 6012
rect 3657 5956 3661 6012
rect 3597 5952 3661 5956
rect 3677 6012 3741 6016
rect 3677 5956 3681 6012
rect 3681 5956 3737 6012
rect 3737 5956 3741 6012
rect 3677 5952 3741 5956
rect 3757 6012 3821 6016
rect 3757 5956 3761 6012
rect 3761 5956 3817 6012
rect 3817 5956 3821 6012
rect 3757 5952 3821 5956
rect 3837 6012 3901 6016
rect 3837 5956 3841 6012
rect 3841 5956 3897 6012
rect 3897 5956 3901 6012
rect 3837 5952 3901 5956
rect 8887 6012 8951 6016
rect 8887 5956 8891 6012
rect 8891 5956 8947 6012
rect 8947 5956 8951 6012
rect 8887 5952 8951 5956
rect 8967 6012 9031 6016
rect 8967 5956 8971 6012
rect 8971 5956 9027 6012
rect 9027 5956 9031 6012
rect 8967 5952 9031 5956
rect 9047 6012 9111 6016
rect 9047 5956 9051 6012
rect 9051 5956 9107 6012
rect 9107 5956 9111 6012
rect 9047 5952 9111 5956
rect 9127 6012 9191 6016
rect 9127 5956 9131 6012
rect 9131 5956 9187 6012
rect 9187 5956 9191 6012
rect 9127 5952 9191 5956
rect 14177 6012 14241 6016
rect 14177 5956 14181 6012
rect 14181 5956 14237 6012
rect 14237 5956 14241 6012
rect 14177 5952 14241 5956
rect 14257 6012 14321 6016
rect 14257 5956 14261 6012
rect 14261 5956 14317 6012
rect 14317 5956 14321 6012
rect 14257 5952 14321 5956
rect 14337 6012 14401 6016
rect 14337 5956 14341 6012
rect 14341 5956 14397 6012
rect 14397 5956 14401 6012
rect 14337 5952 14401 5956
rect 14417 6012 14481 6016
rect 14417 5956 14421 6012
rect 14421 5956 14477 6012
rect 14477 5956 14481 6012
rect 14417 5952 14481 5956
rect 19467 6012 19531 6016
rect 19467 5956 19471 6012
rect 19471 5956 19527 6012
rect 19527 5956 19531 6012
rect 19467 5952 19531 5956
rect 19547 6012 19611 6016
rect 19547 5956 19551 6012
rect 19551 5956 19607 6012
rect 19607 5956 19611 6012
rect 19547 5952 19611 5956
rect 19627 6012 19691 6016
rect 19627 5956 19631 6012
rect 19631 5956 19687 6012
rect 19687 5956 19691 6012
rect 19627 5952 19691 5956
rect 19707 6012 19771 6016
rect 19707 5956 19711 6012
rect 19711 5956 19767 6012
rect 19767 5956 19771 6012
rect 19707 5952 19771 5956
rect 4257 5468 4321 5472
rect 4257 5412 4261 5468
rect 4261 5412 4317 5468
rect 4317 5412 4321 5468
rect 4257 5408 4321 5412
rect 4337 5468 4401 5472
rect 4337 5412 4341 5468
rect 4341 5412 4397 5468
rect 4397 5412 4401 5468
rect 4337 5408 4401 5412
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 9547 5468 9611 5472
rect 9547 5412 9551 5468
rect 9551 5412 9607 5468
rect 9607 5412 9611 5468
rect 9547 5408 9611 5412
rect 9627 5468 9691 5472
rect 9627 5412 9631 5468
rect 9631 5412 9687 5468
rect 9687 5412 9691 5468
rect 9627 5408 9691 5412
rect 9707 5468 9771 5472
rect 9707 5412 9711 5468
rect 9711 5412 9767 5468
rect 9767 5412 9771 5468
rect 9707 5408 9771 5412
rect 9787 5468 9851 5472
rect 9787 5412 9791 5468
rect 9791 5412 9847 5468
rect 9847 5412 9851 5468
rect 9787 5408 9851 5412
rect 14837 5468 14901 5472
rect 14837 5412 14841 5468
rect 14841 5412 14897 5468
rect 14897 5412 14901 5468
rect 14837 5408 14901 5412
rect 14917 5468 14981 5472
rect 14917 5412 14921 5468
rect 14921 5412 14977 5468
rect 14977 5412 14981 5468
rect 14917 5408 14981 5412
rect 14997 5468 15061 5472
rect 14997 5412 15001 5468
rect 15001 5412 15057 5468
rect 15057 5412 15061 5468
rect 14997 5408 15061 5412
rect 15077 5468 15141 5472
rect 15077 5412 15081 5468
rect 15081 5412 15137 5468
rect 15137 5412 15141 5468
rect 15077 5408 15141 5412
rect 20127 5468 20191 5472
rect 20127 5412 20131 5468
rect 20131 5412 20187 5468
rect 20187 5412 20191 5468
rect 20127 5408 20191 5412
rect 20207 5468 20271 5472
rect 20207 5412 20211 5468
rect 20211 5412 20267 5468
rect 20267 5412 20271 5468
rect 20207 5408 20271 5412
rect 20287 5468 20351 5472
rect 20287 5412 20291 5468
rect 20291 5412 20347 5468
rect 20347 5412 20351 5468
rect 20287 5408 20351 5412
rect 20367 5468 20431 5472
rect 20367 5412 20371 5468
rect 20371 5412 20427 5468
rect 20427 5412 20431 5468
rect 20367 5408 20431 5412
rect 3597 4924 3661 4928
rect 3597 4868 3601 4924
rect 3601 4868 3657 4924
rect 3657 4868 3661 4924
rect 3597 4864 3661 4868
rect 3677 4924 3741 4928
rect 3677 4868 3681 4924
rect 3681 4868 3737 4924
rect 3737 4868 3741 4924
rect 3677 4864 3741 4868
rect 3757 4924 3821 4928
rect 3757 4868 3761 4924
rect 3761 4868 3817 4924
rect 3817 4868 3821 4924
rect 3757 4864 3821 4868
rect 3837 4924 3901 4928
rect 3837 4868 3841 4924
rect 3841 4868 3897 4924
rect 3897 4868 3901 4924
rect 3837 4864 3901 4868
rect 8887 4924 8951 4928
rect 8887 4868 8891 4924
rect 8891 4868 8947 4924
rect 8947 4868 8951 4924
rect 8887 4864 8951 4868
rect 8967 4924 9031 4928
rect 8967 4868 8971 4924
rect 8971 4868 9027 4924
rect 9027 4868 9031 4924
rect 8967 4864 9031 4868
rect 9047 4924 9111 4928
rect 9047 4868 9051 4924
rect 9051 4868 9107 4924
rect 9107 4868 9111 4924
rect 9047 4864 9111 4868
rect 9127 4924 9191 4928
rect 9127 4868 9131 4924
rect 9131 4868 9187 4924
rect 9187 4868 9191 4924
rect 9127 4864 9191 4868
rect 14177 4924 14241 4928
rect 14177 4868 14181 4924
rect 14181 4868 14237 4924
rect 14237 4868 14241 4924
rect 14177 4864 14241 4868
rect 14257 4924 14321 4928
rect 14257 4868 14261 4924
rect 14261 4868 14317 4924
rect 14317 4868 14321 4924
rect 14257 4864 14321 4868
rect 14337 4924 14401 4928
rect 14337 4868 14341 4924
rect 14341 4868 14397 4924
rect 14397 4868 14401 4924
rect 14337 4864 14401 4868
rect 14417 4924 14481 4928
rect 14417 4868 14421 4924
rect 14421 4868 14477 4924
rect 14477 4868 14481 4924
rect 14417 4864 14481 4868
rect 19467 4924 19531 4928
rect 19467 4868 19471 4924
rect 19471 4868 19527 4924
rect 19527 4868 19531 4924
rect 19467 4864 19531 4868
rect 19547 4924 19611 4928
rect 19547 4868 19551 4924
rect 19551 4868 19607 4924
rect 19607 4868 19611 4924
rect 19547 4864 19611 4868
rect 19627 4924 19691 4928
rect 19627 4868 19631 4924
rect 19631 4868 19687 4924
rect 19687 4868 19691 4924
rect 19627 4864 19691 4868
rect 19707 4924 19771 4928
rect 19707 4868 19711 4924
rect 19711 4868 19767 4924
rect 19767 4868 19771 4924
rect 19707 4864 19771 4868
rect 4257 4380 4321 4384
rect 4257 4324 4261 4380
rect 4261 4324 4317 4380
rect 4317 4324 4321 4380
rect 4257 4320 4321 4324
rect 4337 4380 4401 4384
rect 4337 4324 4341 4380
rect 4341 4324 4397 4380
rect 4397 4324 4401 4380
rect 4337 4320 4401 4324
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 9547 4380 9611 4384
rect 9547 4324 9551 4380
rect 9551 4324 9607 4380
rect 9607 4324 9611 4380
rect 9547 4320 9611 4324
rect 9627 4380 9691 4384
rect 9627 4324 9631 4380
rect 9631 4324 9687 4380
rect 9687 4324 9691 4380
rect 9627 4320 9691 4324
rect 9707 4380 9771 4384
rect 9707 4324 9711 4380
rect 9711 4324 9767 4380
rect 9767 4324 9771 4380
rect 9707 4320 9771 4324
rect 9787 4380 9851 4384
rect 9787 4324 9791 4380
rect 9791 4324 9847 4380
rect 9847 4324 9851 4380
rect 9787 4320 9851 4324
rect 14837 4380 14901 4384
rect 14837 4324 14841 4380
rect 14841 4324 14897 4380
rect 14897 4324 14901 4380
rect 14837 4320 14901 4324
rect 14917 4380 14981 4384
rect 14917 4324 14921 4380
rect 14921 4324 14977 4380
rect 14977 4324 14981 4380
rect 14917 4320 14981 4324
rect 14997 4380 15061 4384
rect 14997 4324 15001 4380
rect 15001 4324 15057 4380
rect 15057 4324 15061 4380
rect 14997 4320 15061 4324
rect 15077 4380 15141 4384
rect 15077 4324 15081 4380
rect 15081 4324 15137 4380
rect 15137 4324 15141 4380
rect 15077 4320 15141 4324
rect 20127 4380 20191 4384
rect 20127 4324 20131 4380
rect 20131 4324 20187 4380
rect 20187 4324 20191 4380
rect 20127 4320 20191 4324
rect 20207 4380 20271 4384
rect 20207 4324 20211 4380
rect 20211 4324 20267 4380
rect 20267 4324 20271 4380
rect 20207 4320 20271 4324
rect 20287 4380 20351 4384
rect 20287 4324 20291 4380
rect 20291 4324 20347 4380
rect 20347 4324 20351 4380
rect 20287 4320 20351 4324
rect 20367 4380 20431 4384
rect 20367 4324 20371 4380
rect 20371 4324 20427 4380
rect 20427 4324 20431 4380
rect 20367 4320 20431 4324
rect 3597 3836 3661 3840
rect 3597 3780 3601 3836
rect 3601 3780 3657 3836
rect 3657 3780 3661 3836
rect 3597 3776 3661 3780
rect 3677 3836 3741 3840
rect 3677 3780 3681 3836
rect 3681 3780 3737 3836
rect 3737 3780 3741 3836
rect 3677 3776 3741 3780
rect 3757 3836 3821 3840
rect 3757 3780 3761 3836
rect 3761 3780 3817 3836
rect 3817 3780 3821 3836
rect 3757 3776 3821 3780
rect 3837 3836 3901 3840
rect 3837 3780 3841 3836
rect 3841 3780 3897 3836
rect 3897 3780 3901 3836
rect 3837 3776 3901 3780
rect 8887 3836 8951 3840
rect 8887 3780 8891 3836
rect 8891 3780 8947 3836
rect 8947 3780 8951 3836
rect 8887 3776 8951 3780
rect 8967 3836 9031 3840
rect 8967 3780 8971 3836
rect 8971 3780 9027 3836
rect 9027 3780 9031 3836
rect 8967 3776 9031 3780
rect 9047 3836 9111 3840
rect 9047 3780 9051 3836
rect 9051 3780 9107 3836
rect 9107 3780 9111 3836
rect 9047 3776 9111 3780
rect 9127 3836 9191 3840
rect 9127 3780 9131 3836
rect 9131 3780 9187 3836
rect 9187 3780 9191 3836
rect 9127 3776 9191 3780
rect 14177 3836 14241 3840
rect 14177 3780 14181 3836
rect 14181 3780 14237 3836
rect 14237 3780 14241 3836
rect 14177 3776 14241 3780
rect 14257 3836 14321 3840
rect 14257 3780 14261 3836
rect 14261 3780 14317 3836
rect 14317 3780 14321 3836
rect 14257 3776 14321 3780
rect 14337 3836 14401 3840
rect 14337 3780 14341 3836
rect 14341 3780 14397 3836
rect 14397 3780 14401 3836
rect 14337 3776 14401 3780
rect 14417 3836 14481 3840
rect 14417 3780 14421 3836
rect 14421 3780 14477 3836
rect 14477 3780 14481 3836
rect 14417 3776 14481 3780
rect 19467 3836 19531 3840
rect 19467 3780 19471 3836
rect 19471 3780 19527 3836
rect 19527 3780 19531 3836
rect 19467 3776 19531 3780
rect 19547 3836 19611 3840
rect 19547 3780 19551 3836
rect 19551 3780 19607 3836
rect 19607 3780 19611 3836
rect 19547 3776 19611 3780
rect 19627 3836 19691 3840
rect 19627 3780 19631 3836
rect 19631 3780 19687 3836
rect 19687 3780 19691 3836
rect 19627 3776 19691 3780
rect 19707 3836 19771 3840
rect 19707 3780 19711 3836
rect 19711 3780 19767 3836
rect 19767 3780 19771 3836
rect 19707 3776 19771 3780
rect 4257 3292 4321 3296
rect 4257 3236 4261 3292
rect 4261 3236 4317 3292
rect 4317 3236 4321 3292
rect 4257 3232 4321 3236
rect 4337 3292 4401 3296
rect 4337 3236 4341 3292
rect 4341 3236 4397 3292
rect 4397 3236 4401 3292
rect 4337 3232 4401 3236
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 9547 3292 9611 3296
rect 9547 3236 9551 3292
rect 9551 3236 9607 3292
rect 9607 3236 9611 3292
rect 9547 3232 9611 3236
rect 9627 3292 9691 3296
rect 9627 3236 9631 3292
rect 9631 3236 9687 3292
rect 9687 3236 9691 3292
rect 9627 3232 9691 3236
rect 9707 3292 9771 3296
rect 9707 3236 9711 3292
rect 9711 3236 9767 3292
rect 9767 3236 9771 3292
rect 9707 3232 9771 3236
rect 9787 3292 9851 3296
rect 9787 3236 9791 3292
rect 9791 3236 9847 3292
rect 9847 3236 9851 3292
rect 9787 3232 9851 3236
rect 14837 3292 14901 3296
rect 14837 3236 14841 3292
rect 14841 3236 14897 3292
rect 14897 3236 14901 3292
rect 14837 3232 14901 3236
rect 14917 3292 14981 3296
rect 14917 3236 14921 3292
rect 14921 3236 14977 3292
rect 14977 3236 14981 3292
rect 14917 3232 14981 3236
rect 14997 3292 15061 3296
rect 14997 3236 15001 3292
rect 15001 3236 15057 3292
rect 15057 3236 15061 3292
rect 14997 3232 15061 3236
rect 15077 3292 15141 3296
rect 15077 3236 15081 3292
rect 15081 3236 15137 3292
rect 15137 3236 15141 3292
rect 15077 3232 15141 3236
rect 20127 3292 20191 3296
rect 20127 3236 20131 3292
rect 20131 3236 20187 3292
rect 20187 3236 20191 3292
rect 20127 3232 20191 3236
rect 20207 3292 20271 3296
rect 20207 3236 20211 3292
rect 20211 3236 20267 3292
rect 20267 3236 20271 3292
rect 20207 3232 20271 3236
rect 20287 3292 20351 3296
rect 20287 3236 20291 3292
rect 20291 3236 20347 3292
rect 20347 3236 20351 3292
rect 20287 3232 20351 3236
rect 20367 3292 20431 3296
rect 20367 3236 20371 3292
rect 20371 3236 20427 3292
rect 20427 3236 20431 3292
rect 20367 3232 20431 3236
rect 3597 2748 3661 2752
rect 3597 2692 3601 2748
rect 3601 2692 3657 2748
rect 3657 2692 3661 2748
rect 3597 2688 3661 2692
rect 3677 2748 3741 2752
rect 3677 2692 3681 2748
rect 3681 2692 3737 2748
rect 3737 2692 3741 2748
rect 3677 2688 3741 2692
rect 3757 2748 3821 2752
rect 3757 2692 3761 2748
rect 3761 2692 3817 2748
rect 3817 2692 3821 2748
rect 3757 2688 3821 2692
rect 3837 2748 3901 2752
rect 3837 2692 3841 2748
rect 3841 2692 3897 2748
rect 3897 2692 3901 2748
rect 3837 2688 3901 2692
rect 8887 2748 8951 2752
rect 8887 2692 8891 2748
rect 8891 2692 8947 2748
rect 8947 2692 8951 2748
rect 8887 2688 8951 2692
rect 8967 2748 9031 2752
rect 8967 2692 8971 2748
rect 8971 2692 9027 2748
rect 9027 2692 9031 2748
rect 8967 2688 9031 2692
rect 9047 2748 9111 2752
rect 9047 2692 9051 2748
rect 9051 2692 9107 2748
rect 9107 2692 9111 2748
rect 9047 2688 9111 2692
rect 9127 2748 9191 2752
rect 9127 2692 9131 2748
rect 9131 2692 9187 2748
rect 9187 2692 9191 2748
rect 9127 2688 9191 2692
rect 14177 2748 14241 2752
rect 14177 2692 14181 2748
rect 14181 2692 14237 2748
rect 14237 2692 14241 2748
rect 14177 2688 14241 2692
rect 14257 2748 14321 2752
rect 14257 2692 14261 2748
rect 14261 2692 14317 2748
rect 14317 2692 14321 2748
rect 14257 2688 14321 2692
rect 14337 2748 14401 2752
rect 14337 2692 14341 2748
rect 14341 2692 14397 2748
rect 14397 2692 14401 2748
rect 14337 2688 14401 2692
rect 14417 2748 14481 2752
rect 14417 2692 14421 2748
rect 14421 2692 14477 2748
rect 14477 2692 14481 2748
rect 14417 2688 14481 2692
rect 19467 2748 19531 2752
rect 19467 2692 19471 2748
rect 19471 2692 19527 2748
rect 19527 2692 19531 2748
rect 19467 2688 19531 2692
rect 19547 2748 19611 2752
rect 19547 2692 19551 2748
rect 19551 2692 19607 2748
rect 19607 2692 19611 2748
rect 19547 2688 19611 2692
rect 19627 2748 19691 2752
rect 19627 2692 19631 2748
rect 19631 2692 19687 2748
rect 19687 2692 19691 2748
rect 19627 2688 19691 2692
rect 19707 2748 19771 2752
rect 19707 2692 19711 2748
rect 19711 2692 19767 2748
rect 19767 2692 19771 2748
rect 19707 2688 19771 2692
rect 4257 2204 4321 2208
rect 4257 2148 4261 2204
rect 4261 2148 4317 2204
rect 4317 2148 4321 2204
rect 4257 2144 4321 2148
rect 4337 2204 4401 2208
rect 4337 2148 4341 2204
rect 4341 2148 4397 2204
rect 4397 2148 4401 2204
rect 4337 2144 4401 2148
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 9547 2204 9611 2208
rect 9547 2148 9551 2204
rect 9551 2148 9607 2204
rect 9607 2148 9611 2204
rect 9547 2144 9611 2148
rect 9627 2204 9691 2208
rect 9627 2148 9631 2204
rect 9631 2148 9687 2204
rect 9687 2148 9691 2204
rect 9627 2144 9691 2148
rect 9707 2204 9771 2208
rect 9707 2148 9711 2204
rect 9711 2148 9767 2204
rect 9767 2148 9771 2204
rect 9707 2144 9771 2148
rect 9787 2204 9851 2208
rect 9787 2148 9791 2204
rect 9791 2148 9847 2204
rect 9847 2148 9851 2204
rect 9787 2144 9851 2148
rect 14837 2204 14901 2208
rect 14837 2148 14841 2204
rect 14841 2148 14897 2204
rect 14897 2148 14901 2204
rect 14837 2144 14901 2148
rect 14917 2204 14981 2208
rect 14917 2148 14921 2204
rect 14921 2148 14977 2204
rect 14977 2148 14981 2204
rect 14917 2144 14981 2148
rect 14997 2204 15061 2208
rect 14997 2148 15001 2204
rect 15001 2148 15057 2204
rect 15057 2148 15061 2204
rect 14997 2144 15061 2148
rect 15077 2204 15141 2208
rect 15077 2148 15081 2204
rect 15081 2148 15137 2204
rect 15137 2148 15141 2204
rect 15077 2144 15141 2148
rect 20127 2204 20191 2208
rect 20127 2148 20131 2204
rect 20131 2148 20187 2204
rect 20187 2148 20191 2204
rect 20127 2144 20191 2148
rect 20207 2204 20271 2208
rect 20207 2148 20211 2204
rect 20211 2148 20267 2204
rect 20267 2148 20271 2204
rect 20207 2144 20271 2148
rect 20287 2204 20351 2208
rect 20287 2148 20291 2204
rect 20291 2148 20347 2204
rect 20347 2148 20351 2204
rect 20287 2144 20351 2148
rect 20367 2204 20431 2208
rect 20367 2148 20371 2204
rect 20371 2148 20427 2204
rect 20427 2148 20431 2204
rect 20367 2144 20431 2148
<< metal4 >>
rect 3589 22336 3909 22896
rect 3589 22272 3597 22336
rect 3661 22272 3677 22336
rect 3741 22272 3757 22336
rect 3821 22272 3837 22336
rect 3901 22272 3909 22336
rect 3589 21248 3909 22272
rect 3589 21184 3597 21248
rect 3661 21184 3677 21248
rect 3741 21184 3757 21248
rect 3821 21184 3837 21248
rect 3901 21184 3909 21248
rect 3589 20382 3909 21184
rect 3589 20160 3631 20382
rect 3867 20160 3909 20382
rect 3589 20096 3597 20160
rect 3661 20096 3677 20146
rect 3741 20096 3757 20146
rect 3821 20096 3837 20146
rect 3901 20096 3909 20160
rect 3589 19072 3909 20096
rect 3589 19008 3597 19072
rect 3661 19008 3677 19072
rect 3741 19008 3757 19072
rect 3821 19008 3837 19072
rect 3901 19008 3909 19072
rect 3589 17984 3909 19008
rect 3589 17920 3597 17984
rect 3661 17920 3677 17984
rect 3741 17920 3757 17984
rect 3821 17920 3837 17984
rect 3901 17920 3909 17984
rect 3589 16896 3909 17920
rect 3589 16832 3597 16896
rect 3661 16832 3677 16896
rect 3741 16832 3757 16896
rect 3821 16832 3837 16896
rect 3901 16832 3909 16896
rect 3589 15808 3909 16832
rect 3589 15744 3597 15808
rect 3661 15744 3677 15808
rect 3741 15744 3757 15808
rect 3821 15744 3837 15808
rect 3901 15744 3909 15808
rect 3589 15214 3909 15744
rect 3589 14978 3631 15214
rect 3867 14978 3909 15214
rect 3589 14720 3909 14978
rect 3589 14656 3597 14720
rect 3661 14656 3677 14720
rect 3741 14656 3757 14720
rect 3821 14656 3837 14720
rect 3901 14656 3909 14720
rect 3589 13632 3909 14656
rect 3589 13568 3597 13632
rect 3661 13568 3677 13632
rect 3741 13568 3757 13632
rect 3821 13568 3837 13632
rect 3901 13568 3909 13632
rect 3589 12544 3909 13568
rect 3589 12480 3597 12544
rect 3661 12480 3677 12544
rect 3741 12480 3757 12544
rect 3821 12480 3837 12544
rect 3901 12480 3909 12544
rect 3589 11456 3909 12480
rect 3589 11392 3597 11456
rect 3661 11392 3677 11456
rect 3741 11392 3757 11456
rect 3821 11392 3837 11456
rect 3901 11392 3909 11456
rect 3589 10368 3909 11392
rect 3589 10304 3597 10368
rect 3661 10304 3677 10368
rect 3741 10304 3757 10368
rect 3821 10304 3837 10368
rect 3901 10304 3909 10368
rect 3589 10046 3909 10304
rect 3589 9810 3631 10046
rect 3867 9810 3909 10046
rect 3589 9280 3909 9810
rect 3589 9216 3597 9280
rect 3661 9216 3677 9280
rect 3741 9216 3757 9280
rect 3821 9216 3837 9280
rect 3901 9216 3909 9280
rect 3589 8192 3909 9216
rect 3589 8128 3597 8192
rect 3661 8128 3677 8192
rect 3741 8128 3757 8192
rect 3821 8128 3837 8192
rect 3901 8128 3909 8192
rect 3589 7104 3909 8128
rect 3589 7040 3597 7104
rect 3661 7040 3677 7104
rect 3741 7040 3757 7104
rect 3821 7040 3837 7104
rect 3901 7040 3909 7104
rect 3589 6016 3909 7040
rect 3589 5952 3597 6016
rect 3661 5952 3677 6016
rect 3741 5952 3757 6016
rect 3821 5952 3837 6016
rect 3901 5952 3909 6016
rect 3589 4928 3909 5952
rect 3589 4864 3597 4928
rect 3661 4878 3677 4928
rect 3741 4878 3757 4928
rect 3821 4878 3837 4928
rect 3901 4864 3909 4928
rect 3589 4642 3631 4864
rect 3867 4642 3909 4864
rect 3589 3840 3909 4642
rect 3589 3776 3597 3840
rect 3661 3776 3677 3840
rect 3741 3776 3757 3840
rect 3821 3776 3837 3840
rect 3901 3776 3909 3840
rect 3589 2752 3909 3776
rect 3589 2688 3597 2752
rect 3661 2688 3677 2752
rect 3741 2688 3757 2752
rect 3821 2688 3837 2752
rect 3901 2688 3909 2752
rect 3589 2128 3909 2688
rect 4249 22880 4569 22896
rect 4249 22816 4257 22880
rect 4321 22816 4337 22880
rect 4401 22816 4417 22880
rect 4481 22816 4497 22880
rect 4561 22816 4569 22880
rect 4249 21792 4569 22816
rect 4249 21728 4257 21792
rect 4321 21728 4337 21792
rect 4401 21728 4417 21792
rect 4481 21728 4497 21792
rect 4561 21728 4569 21792
rect 4249 21042 4569 21728
rect 4249 20806 4291 21042
rect 4527 20806 4569 21042
rect 4249 20704 4569 20806
rect 4249 20640 4257 20704
rect 4321 20640 4337 20704
rect 4401 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4569 20704
rect 4249 19616 4569 20640
rect 4249 19552 4257 19616
rect 4321 19552 4337 19616
rect 4401 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4569 19616
rect 4249 18528 4569 19552
rect 4249 18464 4257 18528
rect 4321 18464 4337 18528
rect 4401 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4569 18528
rect 4249 17440 4569 18464
rect 4249 17376 4257 17440
rect 4321 17376 4337 17440
rect 4401 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4569 17440
rect 4249 16352 4569 17376
rect 4249 16288 4257 16352
rect 4321 16288 4337 16352
rect 4401 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4569 16352
rect 4249 15874 4569 16288
rect 4249 15638 4291 15874
rect 4527 15638 4569 15874
rect 4249 15264 4569 15638
rect 4249 15200 4257 15264
rect 4321 15200 4337 15264
rect 4401 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4569 15264
rect 4249 14176 4569 15200
rect 4249 14112 4257 14176
rect 4321 14112 4337 14176
rect 4401 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4569 14176
rect 4249 13088 4569 14112
rect 4249 13024 4257 13088
rect 4321 13024 4337 13088
rect 4401 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4569 13088
rect 4249 12000 4569 13024
rect 4249 11936 4257 12000
rect 4321 11936 4337 12000
rect 4401 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4569 12000
rect 4249 10912 4569 11936
rect 4249 10848 4257 10912
rect 4321 10848 4337 10912
rect 4401 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4569 10912
rect 4249 10706 4569 10848
rect 4249 10470 4291 10706
rect 4527 10470 4569 10706
rect 4249 9824 4569 10470
rect 4249 9760 4257 9824
rect 4321 9760 4337 9824
rect 4401 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4569 9824
rect 4249 8736 4569 9760
rect 4249 8672 4257 8736
rect 4321 8672 4337 8736
rect 4401 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4569 8736
rect 4249 7648 4569 8672
rect 4249 7584 4257 7648
rect 4321 7584 4337 7648
rect 4401 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4569 7648
rect 4249 6560 4569 7584
rect 4249 6496 4257 6560
rect 4321 6496 4337 6560
rect 4401 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4569 6560
rect 4249 5538 4569 6496
rect 4249 5472 4291 5538
rect 4527 5472 4569 5538
rect 4249 5408 4257 5472
rect 4561 5408 4569 5472
rect 4249 5302 4291 5408
rect 4527 5302 4569 5408
rect 4249 4384 4569 5302
rect 4249 4320 4257 4384
rect 4321 4320 4337 4384
rect 4401 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4569 4384
rect 4249 3296 4569 4320
rect 4249 3232 4257 3296
rect 4321 3232 4337 3296
rect 4401 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4569 3296
rect 4249 2208 4569 3232
rect 4249 2144 4257 2208
rect 4321 2144 4337 2208
rect 4401 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4569 2208
rect 4249 2128 4569 2144
rect 8879 22336 9199 22896
rect 8879 22272 8887 22336
rect 8951 22272 8967 22336
rect 9031 22272 9047 22336
rect 9111 22272 9127 22336
rect 9191 22272 9199 22336
rect 8879 21248 9199 22272
rect 8879 21184 8887 21248
rect 8951 21184 8967 21248
rect 9031 21184 9047 21248
rect 9111 21184 9127 21248
rect 9191 21184 9199 21248
rect 8879 20382 9199 21184
rect 8879 20160 8921 20382
rect 9157 20160 9199 20382
rect 8879 20096 8887 20160
rect 8951 20096 8967 20146
rect 9031 20096 9047 20146
rect 9111 20096 9127 20146
rect 9191 20096 9199 20160
rect 8879 19072 9199 20096
rect 8879 19008 8887 19072
rect 8951 19008 8967 19072
rect 9031 19008 9047 19072
rect 9111 19008 9127 19072
rect 9191 19008 9199 19072
rect 8879 17984 9199 19008
rect 8879 17920 8887 17984
rect 8951 17920 8967 17984
rect 9031 17920 9047 17984
rect 9111 17920 9127 17984
rect 9191 17920 9199 17984
rect 8879 16896 9199 17920
rect 8879 16832 8887 16896
rect 8951 16832 8967 16896
rect 9031 16832 9047 16896
rect 9111 16832 9127 16896
rect 9191 16832 9199 16896
rect 8879 15808 9199 16832
rect 8879 15744 8887 15808
rect 8951 15744 8967 15808
rect 9031 15744 9047 15808
rect 9111 15744 9127 15808
rect 9191 15744 9199 15808
rect 8879 15214 9199 15744
rect 8879 14978 8921 15214
rect 9157 14978 9199 15214
rect 8879 14720 9199 14978
rect 8879 14656 8887 14720
rect 8951 14656 8967 14720
rect 9031 14656 9047 14720
rect 9111 14656 9127 14720
rect 9191 14656 9199 14720
rect 8879 13632 9199 14656
rect 8879 13568 8887 13632
rect 8951 13568 8967 13632
rect 9031 13568 9047 13632
rect 9111 13568 9127 13632
rect 9191 13568 9199 13632
rect 8879 12544 9199 13568
rect 8879 12480 8887 12544
rect 8951 12480 8967 12544
rect 9031 12480 9047 12544
rect 9111 12480 9127 12544
rect 9191 12480 9199 12544
rect 8879 11456 9199 12480
rect 8879 11392 8887 11456
rect 8951 11392 8967 11456
rect 9031 11392 9047 11456
rect 9111 11392 9127 11456
rect 9191 11392 9199 11456
rect 8879 10368 9199 11392
rect 8879 10304 8887 10368
rect 8951 10304 8967 10368
rect 9031 10304 9047 10368
rect 9111 10304 9127 10368
rect 9191 10304 9199 10368
rect 8879 10046 9199 10304
rect 8879 9810 8921 10046
rect 9157 9810 9199 10046
rect 8879 9280 9199 9810
rect 8879 9216 8887 9280
rect 8951 9216 8967 9280
rect 9031 9216 9047 9280
rect 9111 9216 9127 9280
rect 9191 9216 9199 9280
rect 8879 8192 9199 9216
rect 8879 8128 8887 8192
rect 8951 8128 8967 8192
rect 9031 8128 9047 8192
rect 9111 8128 9127 8192
rect 9191 8128 9199 8192
rect 8879 7104 9199 8128
rect 8879 7040 8887 7104
rect 8951 7040 8967 7104
rect 9031 7040 9047 7104
rect 9111 7040 9127 7104
rect 9191 7040 9199 7104
rect 8879 6016 9199 7040
rect 8879 5952 8887 6016
rect 8951 5952 8967 6016
rect 9031 5952 9047 6016
rect 9111 5952 9127 6016
rect 9191 5952 9199 6016
rect 8879 4928 9199 5952
rect 8879 4864 8887 4928
rect 8951 4878 8967 4928
rect 9031 4878 9047 4928
rect 9111 4878 9127 4928
rect 9191 4864 9199 4928
rect 8879 4642 8921 4864
rect 9157 4642 9199 4864
rect 8879 3840 9199 4642
rect 8879 3776 8887 3840
rect 8951 3776 8967 3840
rect 9031 3776 9047 3840
rect 9111 3776 9127 3840
rect 9191 3776 9199 3840
rect 8879 2752 9199 3776
rect 8879 2688 8887 2752
rect 8951 2688 8967 2752
rect 9031 2688 9047 2752
rect 9111 2688 9127 2752
rect 9191 2688 9199 2752
rect 8879 2128 9199 2688
rect 9539 22880 9859 22896
rect 9539 22816 9547 22880
rect 9611 22816 9627 22880
rect 9691 22816 9707 22880
rect 9771 22816 9787 22880
rect 9851 22816 9859 22880
rect 9539 21792 9859 22816
rect 9539 21728 9547 21792
rect 9611 21728 9627 21792
rect 9691 21728 9707 21792
rect 9771 21728 9787 21792
rect 9851 21728 9859 21792
rect 9539 21042 9859 21728
rect 9539 20806 9581 21042
rect 9817 20806 9859 21042
rect 9539 20704 9859 20806
rect 9539 20640 9547 20704
rect 9611 20640 9627 20704
rect 9691 20640 9707 20704
rect 9771 20640 9787 20704
rect 9851 20640 9859 20704
rect 9539 19616 9859 20640
rect 9539 19552 9547 19616
rect 9611 19552 9627 19616
rect 9691 19552 9707 19616
rect 9771 19552 9787 19616
rect 9851 19552 9859 19616
rect 9539 18528 9859 19552
rect 9539 18464 9547 18528
rect 9611 18464 9627 18528
rect 9691 18464 9707 18528
rect 9771 18464 9787 18528
rect 9851 18464 9859 18528
rect 9539 17440 9859 18464
rect 9539 17376 9547 17440
rect 9611 17376 9627 17440
rect 9691 17376 9707 17440
rect 9771 17376 9787 17440
rect 9851 17376 9859 17440
rect 9539 16352 9859 17376
rect 9539 16288 9547 16352
rect 9611 16288 9627 16352
rect 9691 16288 9707 16352
rect 9771 16288 9787 16352
rect 9851 16288 9859 16352
rect 9539 15874 9859 16288
rect 9539 15638 9581 15874
rect 9817 15638 9859 15874
rect 9539 15264 9859 15638
rect 9539 15200 9547 15264
rect 9611 15200 9627 15264
rect 9691 15200 9707 15264
rect 9771 15200 9787 15264
rect 9851 15200 9859 15264
rect 9539 14176 9859 15200
rect 9539 14112 9547 14176
rect 9611 14112 9627 14176
rect 9691 14112 9707 14176
rect 9771 14112 9787 14176
rect 9851 14112 9859 14176
rect 9539 13088 9859 14112
rect 9539 13024 9547 13088
rect 9611 13024 9627 13088
rect 9691 13024 9707 13088
rect 9771 13024 9787 13088
rect 9851 13024 9859 13088
rect 9539 12000 9859 13024
rect 9539 11936 9547 12000
rect 9611 11936 9627 12000
rect 9691 11936 9707 12000
rect 9771 11936 9787 12000
rect 9851 11936 9859 12000
rect 9539 10912 9859 11936
rect 9539 10848 9547 10912
rect 9611 10848 9627 10912
rect 9691 10848 9707 10912
rect 9771 10848 9787 10912
rect 9851 10848 9859 10912
rect 9539 10706 9859 10848
rect 9539 10470 9581 10706
rect 9817 10470 9859 10706
rect 9539 9824 9859 10470
rect 9539 9760 9547 9824
rect 9611 9760 9627 9824
rect 9691 9760 9707 9824
rect 9771 9760 9787 9824
rect 9851 9760 9859 9824
rect 9539 8736 9859 9760
rect 9539 8672 9547 8736
rect 9611 8672 9627 8736
rect 9691 8672 9707 8736
rect 9771 8672 9787 8736
rect 9851 8672 9859 8736
rect 9539 7648 9859 8672
rect 9539 7584 9547 7648
rect 9611 7584 9627 7648
rect 9691 7584 9707 7648
rect 9771 7584 9787 7648
rect 9851 7584 9859 7648
rect 9539 6560 9859 7584
rect 9539 6496 9547 6560
rect 9611 6496 9627 6560
rect 9691 6496 9707 6560
rect 9771 6496 9787 6560
rect 9851 6496 9859 6560
rect 9539 5538 9859 6496
rect 9539 5472 9581 5538
rect 9817 5472 9859 5538
rect 9539 5408 9547 5472
rect 9851 5408 9859 5472
rect 9539 5302 9581 5408
rect 9817 5302 9859 5408
rect 9539 4384 9859 5302
rect 9539 4320 9547 4384
rect 9611 4320 9627 4384
rect 9691 4320 9707 4384
rect 9771 4320 9787 4384
rect 9851 4320 9859 4384
rect 9539 3296 9859 4320
rect 9539 3232 9547 3296
rect 9611 3232 9627 3296
rect 9691 3232 9707 3296
rect 9771 3232 9787 3296
rect 9851 3232 9859 3296
rect 9539 2208 9859 3232
rect 9539 2144 9547 2208
rect 9611 2144 9627 2208
rect 9691 2144 9707 2208
rect 9771 2144 9787 2208
rect 9851 2144 9859 2208
rect 9539 2128 9859 2144
rect 14169 22336 14489 22896
rect 14169 22272 14177 22336
rect 14241 22272 14257 22336
rect 14321 22272 14337 22336
rect 14401 22272 14417 22336
rect 14481 22272 14489 22336
rect 14169 21248 14489 22272
rect 14169 21184 14177 21248
rect 14241 21184 14257 21248
rect 14321 21184 14337 21248
rect 14401 21184 14417 21248
rect 14481 21184 14489 21248
rect 14169 20382 14489 21184
rect 14169 20160 14211 20382
rect 14447 20160 14489 20382
rect 14169 20096 14177 20160
rect 14241 20096 14257 20146
rect 14321 20096 14337 20146
rect 14401 20096 14417 20146
rect 14481 20096 14489 20160
rect 14169 19072 14489 20096
rect 14169 19008 14177 19072
rect 14241 19008 14257 19072
rect 14321 19008 14337 19072
rect 14401 19008 14417 19072
rect 14481 19008 14489 19072
rect 14169 17984 14489 19008
rect 14169 17920 14177 17984
rect 14241 17920 14257 17984
rect 14321 17920 14337 17984
rect 14401 17920 14417 17984
rect 14481 17920 14489 17984
rect 14169 16896 14489 17920
rect 14169 16832 14177 16896
rect 14241 16832 14257 16896
rect 14321 16832 14337 16896
rect 14401 16832 14417 16896
rect 14481 16832 14489 16896
rect 14169 15808 14489 16832
rect 14169 15744 14177 15808
rect 14241 15744 14257 15808
rect 14321 15744 14337 15808
rect 14401 15744 14417 15808
rect 14481 15744 14489 15808
rect 14169 15214 14489 15744
rect 14169 14978 14211 15214
rect 14447 14978 14489 15214
rect 14169 14720 14489 14978
rect 14169 14656 14177 14720
rect 14241 14656 14257 14720
rect 14321 14656 14337 14720
rect 14401 14656 14417 14720
rect 14481 14656 14489 14720
rect 14169 13632 14489 14656
rect 14169 13568 14177 13632
rect 14241 13568 14257 13632
rect 14321 13568 14337 13632
rect 14401 13568 14417 13632
rect 14481 13568 14489 13632
rect 14169 12544 14489 13568
rect 14169 12480 14177 12544
rect 14241 12480 14257 12544
rect 14321 12480 14337 12544
rect 14401 12480 14417 12544
rect 14481 12480 14489 12544
rect 14169 11456 14489 12480
rect 14169 11392 14177 11456
rect 14241 11392 14257 11456
rect 14321 11392 14337 11456
rect 14401 11392 14417 11456
rect 14481 11392 14489 11456
rect 14169 10368 14489 11392
rect 14169 10304 14177 10368
rect 14241 10304 14257 10368
rect 14321 10304 14337 10368
rect 14401 10304 14417 10368
rect 14481 10304 14489 10368
rect 14169 10046 14489 10304
rect 14169 9810 14211 10046
rect 14447 9810 14489 10046
rect 14169 9280 14489 9810
rect 14169 9216 14177 9280
rect 14241 9216 14257 9280
rect 14321 9216 14337 9280
rect 14401 9216 14417 9280
rect 14481 9216 14489 9280
rect 14169 8192 14489 9216
rect 14169 8128 14177 8192
rect 14241 8128 14257 8192
rect 14321 8128 14337 8192
rect 14401 8128 14417 8192
rect 14481 8128 14489 8192
rect 14169 7104 14489 8128
rect 14169 7040 14177 7104
rect 14241 7040 14257 7104
rect 14321 7040 14337 7104
rect 14401 7040 14417 7104
rect 14481 7040 14489 7104
rect 14169 6016 14489 7040
rect 14169 5952 14177 6016
rect 14241 5952 14257 6016
rect 14321 5952 14337 6016
rect 14401 5952 14417 6016
rect 14481 5952 14489 6016
rect 14169 4928 14489 5952
rect 14169 4864 14177 4928
rect 14241 4878 14257 4928
rect 14321 4878 14337 4928
rect 14401 4878 14417 4928
rect 14481 4864 14489 4928
rect 14169 4642 14211 4864
rect 14447 4642 14489 4864
rect 14169 3840 14489 4642
rect 14169 3776 14177 3840
rect 14241 3776 14257 3840
rect 14321 3776 14337 3840
rect 14401 3776 14417 3840
rect 14481 3776 14489 3840
rect 14169 2752 14489 3776
rect 14169 2688 14177 2752
rect 14241 2688 14257 2752
rect 14321 2688 14337 2752
rect 14401 2688 14417 2752
rect 14481 2688 14489 2752
rect 14169 2128 14489 2688
rect 14829 22880 15149 22896
rect 14829 22816 14837 22880
rect 14901 22816 14917 22880
rect 14981 22816 14997 22880
rect 15061 22816 15077 22880
rect 15141 22816 15149 22880
rect 14829 21792 15149 22816
rect 14829 21728 14837 21792
rect 14901 21728 14917 21792
rect 14981 21728 14997 21792
rect 15061 21728 15077 21792
rect 15141 21728 15149 21792
rect 14829 21042 15149 21728
rect 14829 20806 14871 21042
rect 15107 20806 15149 21042
rect 14829 20704 15149 20806
rect 14829 20640 14837 20704
rect 14901 20640 14917 20704
rect 14981 20640 14997 20704
rect 15061 20640 15077 20704
rect 15141 20640 15149 20704
rect 14829 19616 15149 20640
rect 14829 19552 14837 19616
rect 14901 19552 14917 19616
rect 14981 19552 14997 19616
rect 15061 19552 15077 19616
rect 15141 19552 15149 19616
rect 14829 18528 15149 19552
rect 14829 18464 14837 18528
rect 14901 18464 14917 18528
rect 14981 18464 14997 18528
rect 15061 18464 15077 18528
rect 15141 18464 15149 18528
rect 14829 17440 15149 18464
rect 14829 17376 14837 17440
rect 14901 17376 14917 17440
rect 14981 17376 14997 17440
rect 15061 17376 15077 17440
rect 15141 17376 15149 17440
rect 14829 16352 15149 17376
rect 14829 16288 14837 16352
rect 14901 16288 14917 16352
rect 14981 16288 14997 16352
rect 15061 16288 15077 16352
rect 15141 16288 15149 16352
rect 14829 15874 15149 16288
rect 14829 15638 14871 15874
rect 15107 15638 15149 15874
rect 14829 15264 15149 15638
rect 14829 15200 14837 15264
rect 14901 15200 14917 15264
rect 14981 15200 14997 15264
rect 15061 15200 15077 15264
rect 15141 15200 15149 15264
rect 14829 14176 15149 15200
rect 14829 14112 14837 14176
rect 14901 14112 14917 14176
rect 14981 14112 14997 14176
rect 15061 14112 15077 14176
rect 15141 14112 15149 14176
rect 14829 13088 15149 14112
rect 14829 13024 14837 13088
rect 14901 13024 14917 13088
rect 14981 13024 14997 13088
rect 15061 13024 15077 13088
rect 15141 13024 15149 13088
rect 14829 12000 15149 13024
rect 14829 11936 14837 12000
rect 14901 11936 14917 12000
rect 14981 11936 14997 12000
rect 15061 11936 15077 12000
rect 15141 11936 15149 12000
rect 14829 10912 15149 11936
rect 14829 10848 14837 10912
rect 14901 10848 14917 10912
rect 14981 10848 14997 10912
rect 15061 10848 15077 10912
rect 15141 10848 15149 10912
rect 14829 10706 15149 10848
rect 14829 10470 14871 10706
rect 15107 10470 15149 10706
rect 14829 9824 15149 10470
rect 14829 9760 14837 9824
rect 14901 9760 14917 9824
rect 14981 9760 14997 9824
rect 15061 9760 15077 9824
rect 15141 9760 15149 9824
rect 14829 8736 15149 9760
rect 14829 8672 14837 8736
rect 14901 8672 14917 8736
rect 14981 8672 14997 8736
rect 15061 8672 15077 8736
rect 15141 8672 15149 8736
rect 14829 7648 15149 8672
rect 14829 7584 14837 7648
rect 14901 7584 14917 7648
rect 14981 7584 14997 7648
rect 15061 7584 15077 7648
rect 15141 7584 15149 7648
rect 14829 6560 15149 7584
rect 14829 6496 14837 6560
rect 14901 6496 14917 6560
rect 14981 6496 14997 6560
rect 15061 6496 15077 6560
rect 15141 6496 15149 6560
rect 14829 5538 15149 6496
rect 14829 5472 14871 5538
rect 15107 5472 15149 5538
rect 14829 5408 14837 5472
rect 15141 5408 15149 5472
rect 14829 5302 14871 5408
rect 15107 5302 15149 5408
rect 14829 4384 15149 5302
rect 14829 4320 14837 4384
rect 14901 4320 14917 4384
rect 14981 4320 14997 4384
rect 15061 4320 15077 4384
rect 15141 4320 15149 4384
rect 14829 3296 15149 4320
rect 14829 3232 14837 3296
rect 14901 3232 14917 3296
rect 14981 3232 14997 3296
rect 15061 3232 15077 3296
rect 15141 3232 15149 3296
rect 14829 2208 15149 3232
rect 14829 2144 14837 2208
rect 14901 2144 14917 2208
rect 14981 2144 14997 2208
rect 15061 2144 15077 2208
rect 15141 2144 15149 2208
rect 14829 2128 15149 2144
rect 19459 22336 19779 22896
rect 19459 22272 19467 22336
rect 19531 22272 19547 22336
rect 19611 22272 19627 22336
rect 19691 22272 19707 22336
rect 19771 22272 19779 22336
rect 19459 21248 19779 22272
rect 19459 21184 19467 21248
rect 19531 21184 19547 21248
rect 19611 21184 19627 21248
rect 19691 21184 19707 21248
rect 19771 21184 19779 21248
rect 19459 20382 19779 21184
rect 19459 20160 19501 20382
rect 19737 20160 19779 20382
rect 19459 20096 19467 20160
rect 19531 20096 19547 20146
rect 19611 20096 19627 20146
rect 19691 20096 19707 20146
rect 19771 20096 19779 20160
rect 19459 19072 19779 20096
rect 19459 19008 19467 19072
rect 19531 19008 19547 19072
rect 19611 19008 19627 19072
rect 19691 19008 19707 19072
rect 19771 19008 19779 19072
rect 19459 17984 19779 19008
rect 19459 17920 19467 17984
rect 19531 17920 19547 17984
rect 19611 17920 19627 17984
rect 19691 17920 19707 17984
rect 19771 17920 19779 17984
rect 19459 16896 19779 17920
rect 19459 16832 19467 16896
rect 19531 16832 19547 16896
rect 19611 16832 19627 16896
rect 19691 16832 19707 16896
rect 19771 16832 19779 16896
rect 19459 15808 19779 16832
rect 19459 15744 19467 15808
rect 19531 15744 19547 15808
rect 19611 15744 19627 15808
rect 19691 15744 19707 15808
rect 19771 15744 19779 15808
rect 19459 15214 19779 15744
rect 19459 14978 19501 15214
rect 19737 14978 19779 15214
rect 19459 14720 19779 14978
rect 19459 14656 19467 14720
rect 19531 14656 19547 14720
rect 19611 14656 19627 14720
rect 19691 14656 19707 14720
rect 19771 14656 19779 14720
rect 19459 13632 19779 14656
rect 19459 13568 19467 13632
rect 19531 13568 19547 13632
rect 19611 13568 19627 13632
rect 19691 13568 19707 13632
rect 19771 13568 19779 13632
rect 19459 12544 19779 13568
rect 19459 12480 19467 12544
rect 19531 12480 19547 12544
rect 19611 12480 19627 12544
rect 19691 12480 19707 12544
rect 19771 12480 19779 12544
rect 19459 11456 19779 12480
rect 19459 11392 19467 11456
rect 19531 11392 19547 11456
rect 19611 11392 19627 11456
rect 19691 11392 19707 11456
rect 19771 11392 19779 11456
rect 19459 10368 19779 11392
rect 19459 10304 19467 10368
rect 19531 10304 19547 10368
rect 19611 10304 19627 10368
rect 19691 10304 19707 10368
rect 19771 10304 19779 10368
rect 19459 10046 19779 10304
rect 19459 9810 19501 10046
rect 19737 9810 19779 10046
rect 19459 9280 19779 9810
rect 19459 9216 19467 9280
rect 19531 9216 19547 9280
rect 19611 9216 19627 9280
rect 19691 9216 19707 9280
rect 19771 9216 19779 9280
rect 19459 8192 19779 9216
rect 19459 8128 19467 8192
rect 19531 8128 19547 8192
rect 19611 8128 19627 8192
rect 19691 8128 19707 8192
rect 19771 8128 19779 8192
rect 19459 7104 19779 8128
rect 19459 7040 19467 7104
rect 19531 7040 19547 7104
rect 19611 7040 19627 7104
rect 19691 7040 19707 7104
rect 19771 7040 19779 7104
rect 19459 6016 19779 7040
rect 19459 5952 19467 6016
rect 19531 5952 19547 6016
rect 19611 5952 19627 6016
rect 19691 5952 19707 6016
rect 19771 5952 19779 6016
rect 19459 4928 19779 5952
rect 19459 4864 19467 4928
rect 19531 4878 19547 4928
rect 19611 4878 19627 4928
rect 19691 4878 19707 4928
rect 19771 4864 19779 4928
rect 19459 4642 19501 4864
rect 19737 4642 19779 4864
rect 19459 3840 19779 4642
rect 19459 3776 19467 3840
rect 19531 3776 19547 3840
rect 19611 3776 19627 3840
rect 19691 3776 19707 3840
rect 19771 3776 19779 3840
rect 19459 2752 19779 3776
rect 19459 2688 19467 2752
rect 19531 2688 19547 2752
rect 19611 2688 19627 2752
rect 19691 2688 19707 2752
rect 19771 2688 19779 2752
rect 19459 2128 19779 2688
rect 20119 22880 20439 22896
rect 20119 22816 20127 22880
rect 20191 22816 20207 22880
rect 20271 22816 20287 22880
rect 20351 22816 20367 22880
rect 20431 22816 20439 22880
rect 20119 21792 20439 22816
rect 20119 21728 20127 21792
rect 20191 21728 20207 21792
rect 20271 21728 20287 21792
rect 20351 21728 20367 21792
rect 20431 21728 20439 21792
rect 20119 21042 20439 21728
rect 20119 20806 20161 21042
rect 20397 20806 20439 21042
rect 20119 20704 20439 20806
rect 20119 20640 20127 20704
rect 20191 20640 20207 20704
rect 20271 20640 20287 20704
rect 20351 20640 20367 20704
rect 20431 20640 20439 20704
rect 20119 19616 20439 20640
rect 20119 19552 20127 19616
rect 20191 19552 20207 19616
rect 20271 19552 20287 19616
rect 20351 19552 20367 19616
rect 20431 19552 20439 19616
rect 20119 18528 20439 19552
rect 20119 18464 20127 18528
rect 20191 18464 20207 18528
rect 20271 18464 20287 18528
rect 20351 18464 20367 18528
rect 20431 18464 20439 18528
rect 20119 17440 20439 18464
rect 20119 17376 20127 17440
rect 20191 17376 20207 17440
rect 20271 17376 20287 17440
rect 20351 17376 20367 17440
rect 20431 17376 20439 17440
rect 20119 16352 20439 17376
rect 20119 16288 20127 16352
rect 20191 16288 20207 16352
rect 20271 16288 20287 16352
rect 20351 16288 20367 16352
rect 20431 16288 20439 16352
rect 20119 15874 20439 16288
rect 20119 15638 20161 15874
rect 20397 15638 20439 15874
rect 20119 15264 20439 15638
rect 20119 15200 20127 15264
rect 20191 15200 20207 15264
rect 20271 15200 20287 15264
rect 20351 15200 20367 15264
rect 20431 15200 20439 15264
rect 20119 14176 20439 15200
rect 20119 14112 20127 14176
rect 20191 14112 20207 14176
rect 20271 14112 20287 14176
rect 20351 14112 20367 14176
rect 20431 14112 20439 14176
rect 20119 13088 20439 14112
rect 20119 13024 20127 13088
rect 20191 13024 20207 13088
rect 20271 13024 20287 13088
rect 20351 13024 20367 13088
rect 20431 13024 20439 13088
rect 20119 12000 20439 13024
rect 20119 11936 20127 12000
rect 20191 11936 20207 12000
rect 20271 11936 20287 12000
rect 20351 11936 20367 12000
rect 20431 11936 20439 12000
rect 20119 10912 20439 11936
rect 20119 10848 20127 10912
rect 20191 10848 20207 10912
rect 20271 10848 20287 10912
rect 20351 10848 20367 10912
rect 20431 10848 20439 10912
rect 20119 10706 20439 10848
rect 20119 10470 20161 10706
rect 20397 10470 20439 10706
rect 20119 9824 20439 10470
rect 20119 9760 20127 9824
rect 20191 9760 20207 9824
rect 20271 9760 20287 9824
rect 20351 9760 20367 9824
rect 20431 9760 20439 9824
rect 20119 8736 20439 9760
rect 20119 8672 20127 8736
rect 20191 8672 20207 8736
rect 20271 8672 20287 8736
rect 20351 8672 20367 8736
rect 20431 8672 20439 8736
rect 20119 7648 20439 8672
rect 20119 7584 20127 7648
rect 20191 7584 20207 7648
rect 20271 7584 20287 7648
rect 20351 7584 20367 7648
rect 20431 7584 20439 7648
rect 20119 6560 20439 7584
rect 20119 6496 20127 6560
rect 20191 6496 20207 6560
rect 20271 6496 20287 6560
rect 20351 6496 20367 6560
rect 20431 6496 20439 6560
rect 20119 5538 20439 6496
rect 20119 5472 20161 5538
rect 20397 5472 20439 5538
rect 20119 5408 20127 5472
rect 20431 5408 20439 5472
rect 20119 5302 20161 5408
rect 20397 5302 20439 5408
rect 20119 4384 20439 5302
rect 20119 4320 20127 4384
rect 20191 4320 20207 4384
rect 20271 4320 20287 4384
rect 20351 4320 20367 4384
rect 20431 4320 20439 4384
rect 20119 3296 20439 4320
rect 20119 3232 20127 3296
rect 20191 3232 20207 3296
rect 20271 3232 20287 3296
rect 20351 3232 20367 3296
rect 20431 3232 20439 3296
rect 20119 2208 20439 3232
rect 20119 2144 20127 2208
rect 20191 2144 20207 2208
rect 20271 2144 20287 2208
rect 20351 2144 20367 2208
rect 20431 2144 20439 2208
rect 20119 2128 20439 2144
<< via4 >>
rect 3631 20160 3867 20382
rect 3631 20146 3661 20160
rect 3661 20146 3677 20160
rect 3677 20146 3741 20160
rect 3741 20146 3757 20160
rect 3757 20146 3821 20160
rect 3821 20146 3837 20160
rect 3837 20146 3867 20160
rect 3631 14978 3867 15214
rect 3631 9810 3867 10046
rect 3631 4864 3661 4878
rect 3661 4864 3677 4878
rect 3677 4864 3741 4878
rect 3741 4864 3757 4878
rect 3757 4864 3821 4878
rect 3821 4864 3837 4878
rect 3837 4864 3867 4878
rect 3631 4642 3867 4864
rect 4291 20806 4527 21042
rect 4291 15638 4527 15874
rect 4291 10470 4527 10706
rect 4291 5472 4527 5538
rect 4291 5408 4321 5472
rect 4321 5408 4337 5472
rect 4337 5408 4401 5472
rect 4401 5408 4417 5472
rect 4417 5408 4481 5472
rect 4481 5408 4497 5472
rect 4497 5408 4527 5472
rect 4291 5302 4527 5408
rect 8921 20160 9157 20382
rect 8921 20146 8951 20160
rect 8951 20146 8967 20160
rect 8967 20146 9031 20160
rect 9031 20146 9047 20160
rect 9047 20146 9111 20160
rect 9111 20146 9127 20160
rect 9127 20146 9157 20160
rect 8921 14978 9157 15214
rect 8921 9810 9157 10046
rect 8921 4864 8951 4878
rect 8951 4864 8967 4878
rect 8967 4864 9031 4878
rect 9031 4864 9047 4878
rect 9047 4864 9111 4878
rect 9111 4864 9127 4878
rect 9127 4864 9157 4878
rect 8921 4642 9157 4864
rect 9581 20806 9817 21042
rect 9581 15638 9817 15874
rect 9581 10470 9817 10706
rect 9581 5472 9817 5538
rect 9581 5408 9611 5472
rect 9611 5408 9627 5472
rect 9627 5408 9691 5472
rect 9691 5408 9707 5472
rect 9707 5408 9771 5472
rect 9771 5408 9787 5472
rect 9787 5408 9817 5472
rect 9581 5302 9817 5408
rect 14211 20160 14447 20382
rect 14211 20146 14241 20160
rect 14241 20146 14257 20160
rect 14257 20146 14321 20160
rect 14321 20146 14337 20160
rect 14337 20146 14401 20160
rect 14401 20146 14417 20160
rect 14417 20146 14447 20160
rect 14211 14978 14447 15214
rect 14211 9810 14447 10046
rect 14211 4864 14241 4878
rect 14241 4864 14257 4878
rect 14257 4864 14321 4878
rect 14321 4864 14337 4878
rect 14337 4864 14401 4878
rect 14401 4864 14417 4878
rect 14417 4864 14447 4878
rect 14211 4642 14447 4864
rect 14871 20806 15107 21042
rect 14871 15638 15107 15874
rect 14871 10470 15107 10706
rect 14871 5472 15107 5538
rect 14871 5408 14901 5472
rect 14901 5408 14917 5472
rect 14917 5408 14981 5472
rect 14981 5408 14997 5472
rect 14997 5408 15061 5472
rect 15061 5408 15077 5472
rect 15077 5408 15107 5472
rect 14871 5302 15107 5408
rect 19501 20160 19737 20382
rect 19501 20146 19531 20160
rect 19531 20146 19547 20160
rect 19547 20146 19611 20160
rect 19611 20146 19627 20160
rect 19627 20146 19691 20160
rect 19691 20146 19707 20160
rect 19707 20146 19737 20160
rect 19501 14978 19737 15214
rect 19501 9810 19737 10046
rect 19501 4864 19531 4878
rect 19531 4864 19547 4878
rect 19547 4864 19611 4878
rect 19611 4864 19627 4878
rect 19627 4864 19691 4878
rect 19691 4864 19707 4878
rect 19707 4864 19737 4878
rect 19501 4642 19737 4864
rect 20161 20806 20397 21042
rect 20161 15638 20397 15874
rect 20161 10470 20397 10706
rect 20161 5472 20397 5538
rect 20161 5408 20191 5472
rect 20191 5408 20207 5472
rect 20207 5408 20271 5472
rect 20271 5408 20287 5472
rect 20287 5408 20351 5472
rect 20351 5408 20367 5472
rect 20367 5408 20397 5472
rect 20161 5302 20397 5408
<< metal5 >>
rect 1056 21042 22312 21084
rect 1056 20806 4291 21042
rect 4527 20806 9581 21042
rect 9817 20806 14871 21042
rect 15107 20806 20161 21042
rect 20397 20806 22312 21042
rect 1056 20764 22312 20806
rect 1056 20382 22312 20424
rect 1056 20146 3631 20382
rect 3867 20146 8921 20382
rect 9157 20146 14211 20382
rect 14447 20146 19501 20382
rect 19737 20146 22312 20382
rect 1056 20104 22312 20146
rect 1056 15874 22312 15916
rect 1056 15638 4291 15874
rect 4527 15638 9581 15874
rect 9817 15638 14871 15874
rect 15107 15638 20161 15874
rect 20397 15638 22312 15874
rect 1056 15596 22312 15638
rect 1056 15214 22312 15256
rect 1056 14978 3631 15214
rect 3867 14978 8921 15214
rect 9157 14978 14211 15214
rect 14447 14978 19501 15214
rect 19737 14978 22312 15214
rect 1056 14936 22312 14978
rect 1056 10706 22312 10748
rect 1056 10470 4291 10706
rect 4527 10470 9581 10706
rect 9817 10470 14871 10706
rect 15107 10470 20161 10706
rect 20397 10470 22312 10706
rect 1056 10428 22312 10470
rect 1056 10046 22312 10088
rect 1056 9810 3631 10046
rect 3867 9810 8921 10046
rect 9157 9810 14211 10046
rect 14447 9810 19501 10046
rect 19737 9810 22312 10046
rect 1056 9768 22312 9810
rect 1056 5538 22312 5580
rect 1056 5302 4291 5538
rect 4527 5302 9581 5538
rect 9817 5302 14871 5538
rect 15107 5302 20161 5538
rect 20397 5302 22312 5538
rect 1056 5260 22312 5302
rect 1056 4878 22312 4920
rect 1056 4642 3631 4878
rect 3867 4642 8921 4878
rect 9157 4642 14211 4878
rect 14447 4642 19501 4878
rect 19737 4642 22312 4878
rect 1056 4600 22312 4642
use sky130_fd_sc_hd__and4_1  _442_
timestamp 0
transform -1 0 18032 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _443_
timestamp 0
transform 1 0 15916 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _444_
timestamp 0
transform -1 0 17112 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _445_
timestamp 0
transform 1 0 16192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _446_
timestamp 0
transform -1 0 17756 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _447_
timestamp 0
transform -1 0 20148 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _448_
timestamp 0
transform -1 0 19688 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _449_
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _450_
timestamp 0
transform 1 0 18216 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _451_
timestamp 0
transform -1 0 20240 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _452_
timestamp 0
transform -1 0 19780 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _453_
timestamp 0
transform -1 0 19044 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _454_
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _455_
timestamp 0
transform -1 0 15732 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _456_
timestamp 0
transform -1 0 14720 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _457_
timestamp 0
transform 1 0 14260 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _458_
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _459_
timestamp 0
transform 1 0 6348 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _460_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _461_
timestamp 0
transform -1 0 8096 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _462_
timestamp 0
transform 1 0 19780 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _463_
timestamp 0
transform -1 0 21068 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _464_
timestamp 0
transform 1 0 20424 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _465_
timestamp 0
transform 1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 0
transform -1 0 10672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _467_
timestamp 0
transform 1 0 6624 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 0
transform -1 0 8464 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 0
transform -1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 0
transform -1 0 7360 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp 0
transform 1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 0
transform -1 0 12880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _473_
timestamp 0
transform 1 0 6440 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 0
transform -1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _475_
timestamp 0
transform -1 0 7728 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _476_
timestamp 0
transform -1 0 7728 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _477_
timestamp 0
transform -1 0 8556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _478_
timestamp 0
transform 1 0 6532 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _479_
timestamp 0
transform 1 0 6992 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _480_
timestamp 0
transform -1 0 7728 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _481_
timestamp 0
transform 1 0 7268 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _482_
timestamp 0
transform 1 0 7820 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _483_
timestamp 0
transform -1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _484_
timestamp 0
transform -1 0 6716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _485_
timestamp 0
transform 1 0 3404 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _486_
timestamp 0
transform -1 0 4876 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _487_
timestamp 0
transform -1 0 5060 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _488_
timestamp 0
transform -1 0 5704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _489_
timestamp 0
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _490_
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _491_
timestamp 0
transform 1 0 5336 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _492_
timestamp 0
transform -1 0 5336 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _493_
timestamp 0
transform -1 0 4784 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _494_
timestamp 0
transform 1 0 4416 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _495_
timestamp 0
transform 1 0 4508 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _496_
timestamp 0
transform -1 0 4692 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _497_
timestamp 0
transform -1 0 4784 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _498_
timestamp 0
transform -1 0 5060 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _499_
timestamp 0
transform -1 0 4600 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _500_
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _501_
timestamp 0
transform 1 0 2300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _502_
timestamp 0
transform 1 0 13248 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _503_
timestamp 0
transform 1 0 13248 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _504_
timestamp 0
transform 1 0 12420 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _505_
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _506_
timestamp 0
transform 1 0 12236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _507_
timestamp 0
transform 1 0 13248 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _508_
timestamp 0
transform 1 0 12972 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _509_
timestamp 0
transform 1 0 12236 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _510_
timestamp 0
transform 1 0 12880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _511_
timestamp 0
transform 1 0 12880 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _512_
timestamp 0
transform -1 0 13064 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _513_
timestamp 0
transform 1 0 12420 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _514_
timestamp 0
transform 1 0 12512 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _515_
timestamp 0
transform 1 0 12880 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _516_
timestamp 0
transform 1 0 12696 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _517_
timestamp 0
transform 1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _518_
timestamp 0
transform 1 0 13156 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _519_
timestamp 0
transform 1 0 13248 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _520_
timestamp 0
transform -1 0 17940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _521_
timestamp 0
transform -1 0 16836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _522_
timestamp 0
transform -1 0 16192 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _523_
timestamp 0
transform 1 0 17756 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _524_
timestamp 0
transform -1 0 20148 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _525_
timestamp 0
transform -1 0 18492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _526_
timestamp 0
transform 1 0 18216 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _527_
timestamp 0
transform -1 0 20332 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _528_
timestamp 0
transform -1 0 19780 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _529_
timestamp 0
transform 1 0 13064 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _530_
timestamp 0
transform -1 0 15272 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _531_
timestamp 0
transform -1 0 13616 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _532_
timestamp 0
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _533_
timestamp 0
transform 1 0 6532 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _534_
timestamp 0
transform -1 0 7636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _535_
timestamp 0
transform -1 0 19780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _536_
timestamp 0
transform -1 0 21252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _537_
timestamp 0
transform -1 0 21068 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _538_
timestamp 0
transform -1 0 15272 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _539_
timestamp 0
transform 1 0 9752 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _540_
timestamp 0
transform -1 0 15824 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _541_
timestamp 0
transform -1 0 12052 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _542_
timestamp 0
transform 1 0 12512 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _543_
timestamp 0
transform -1 0 12512 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _544_
timestamp 0
transform -1 0 10396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _545_
timestamp 0
transform -1 0 9844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _546_
timestamp 0
transform -1 0 11316 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _547_
timestamp 0
transform 1 0 15824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _548_
timestamp 0
transform 1 0 8924 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _549_
timestamp 0
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _550_
timestamp 0
transform -1 0 11408 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _551_
timestamp 0
transform 1 0 9292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _552_
timestamp 0
transform -1 0 12420 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _553_
timestamp 0
transform -1 0 10580 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _554_
timestamp 0
transform 1 0 9936 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _555_
timestamp 0
transform -1 0 11224 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _556_
timestamp 0
transform -1 0 9752 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _557_
timestamp 0
transform 1 0 10212 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _558_
timestamp 0
transform -1 0 12420 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _559_
timestamp 0
transform -1 0 11224 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _560_
timestamp 0
transform 1 0 10396 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _561_
timestamp 0
transform -1 0 12328 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _562_
timestamp 0
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _563_
timestamp 0
transform 1 0 13248 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _564_
timestamp 0
transform 1 0 14812 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _565_
timestamp 0
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _566_
timestamp 0
transform -1 0 14260 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 0
transform -1 0 13524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _568_
timestamp 0
transform -1 0 13892 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 0
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _570_
timestamp 0
transform -1 0 17848 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 0
transform -1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _572_
timestamp 0
transform 1 0 16928 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 0
transform -1 0 18952 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _574_
timestamp 0
transform -1 0 18032 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp 0
transform -1 0 17020 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _576_
timestamp 0
transform -1 0 19136 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _577_
timestamp 0
transform -1 0 18768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _578_
timestamp 0
transform 1 0 19964 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _579_
timestamp 0
transform -1 0 20240 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _580_
timestamp 0
transform 1 0 18400 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _581_
timestamp 0
transform -1 0 19136 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _582_
timestamp 0
transform 1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _583_
timestamp 0
transform 1 0 19780 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _584_
timestamp 0
transform -1 0 20516 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _585_
timestamp 0
transform -1 0 21712 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _586_
timestamp 0
transform 1 0 21068 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _587_
timestamp 0
transform -1 0 20424 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _588_
timestamp 0
transform -1 0 19136 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _589_
timestamp 0
transform 1 0 18584 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _590_
timestamp 0
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _591_
timestamp 0
transform -1 0 18216 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _592_
timestamp 0
transform -1 0 17572 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _593_
timestamp 0
transform -1 0 20976 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _594_
timestamp 0
transform -1 0 19780 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _595_
timestamp 0
transform 1 0 20148 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _596_
timestamp 0
transform 1 0 20240 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _597_
timestamp 0
transform 1 0 14076 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _598_
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _599_
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _600_
timestamp 0
transform -1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _601_
timestamp 0
transform -1 0 12328 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _602_
timestamp 0
transform -1 0 13708 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _603_
timestamp 0
transform 1 0 11592 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _604_
timestamp 0
transform -1 0 12420 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _605_
timestamp 0
transform -1 0 11960 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _606_
timestamp 0
transform 1 0 10672 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _607_
timestamp 0
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _608_
timestamp 0
transform -1 0 12144 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _609_
timestamp 0
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _610_
timestamp 0
transform -1 0 11868 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _611_
timestamp 0
transform -1 0 11868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _612_
timestamp 0
transform -1 0 13984 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _613_
timestamp 0
transform 1 0 13800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _614_
timestamp 0
transform 1 0 12052 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _615_
timestamp 0
transform 1 0 11868 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _616_
timestamp 0
transform -1 0 9936 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _617_
timestamp 0
transform -1 0 10672 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _618_
timestamp 0
transform 1 0 9660 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _619_
timestamp 0
transform -1 0 10212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _620_
timestamp 0
transform 1 0 9844 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _621_
timestamp 0
transform -1 0 9476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _622_
timestamp 0
transform 1 0 7360 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _623_
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _624_
timestamp 0
transform 1 0 8004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _625_
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _626_
timestamp 0
transform 1 0 7544 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _627_
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_2  _628_
timestamp 0
transform 1 0 8648 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _629_
timestamp 0
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _630_
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _631_
timestamp 0
transform 1 0 8004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _632_
timestamp 0
transform 1 0 8188 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _633_
timestamp 0
transform 1 0 9292 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _634_
timestamp 0
transform 1 0 9384 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _635_
timestamp 0
transform 1 0 8832 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _636_
timestamp 0
transform 1 0 9016 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _637_
timestamp 0
transform -1 0 10856 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _638_
timestamp 0
transform -1 0 10488 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _639_
timestamp 0
transform -1 0 11960 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _640_
timestamp 0
transform -1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _641_
timestamp 0
transform -1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_4  _642_
timestamp 0
transform 1 0 9844 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__o22ai_1  _643_
timestamp 0
transform 1 0 10948 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _644_
timestamp 0
transform 1 0 12420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _645_
timestamp 0
transform 1 0 10948 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _646_
timestamp 0
transform -1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _647_
timestamp 0
transform -1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _648_
timestamp 0
transform 1 0 11776 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _649_
timestamp 0
transform 1 0 9108 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _650_
timestamp 0
transform 1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _651_
timestamp 0
transform 1 0 9752 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _652_
timestamp 0
transform 1 0 10304 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a311oi_1  _653_
timestamp 0
transform 1 0 9568 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _654_
timestamp 0
transform 1 0 15088 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _655_
timestamp 0
transform 1 0 15364 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _656_
timestamp 0
transform 1 0 15824 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _657_
timestamp 0
transform -1 0 16560 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _658_
timestamp 0
transform -1 0 21620 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _659_
timestamp 0
transform -1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _660_
timestamp 0
transform 1 0 20516 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _661_
timestamp 0
transform 1 0 21620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _662_
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _663_
timestamp 0
transform 1 0 20056 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _664_
timestamp 0
transform 1 0 20240 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _665_
timestamp 0
transform 1 0 18308 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _666_
timestamp 0
transform 1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _667_
timestamp 0
transform -1 0 17480 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _668_
timestamp 0
transform -1 0 16560 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _669_
timestamp 0
transform -1 0 17112 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _670_
timestamp 0
transform -1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _671_
timestamp 0
transform -1 0 16560 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _672_
timestamp 0
transform -1 0 16100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _673_
timestamp 0
transform 1 0 12972 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _674_
timestamp 0
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _675_
timestamp 0
transform 1 0 20240 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _676_
timestamp 0
transform -1 0 20976 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _677_
timestamp 0
transform -1 0 20976 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _678_
timestamp 0
transform -1 0 20240 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _679_
timestamp 0
transform 1 0 19320 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _680_
timestamp 0
transform -1 0 19964 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _681_
timestamp 0
transform -1 0 19136 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _682_
timestamp 0
transform -1 0 17940 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _683_
timestamp 0
transform -1 0 19688 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _684_
timestamp 0
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _685_
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _686_
timestamp 0
transform 1 0 17112 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _687_
timestamp 0
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _688_
timestamp 0
transform 1 0 16560 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _689_
timestamp 0
transform 1 0 17572 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _690_
timestamp 0
transform -1 0 19688 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _691_
timestamp 0
transform -1 0 19412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _692_
timestamp 0
transform -1 0 14536 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _693_
timestamp 0
transform -1 0 13984 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _694_
timestamp 0
transform 1 0 10488 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _695_
timestamp 0
transform 1 0 9660 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _696_
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _697_
timestamp 0
transform 1 0 9476 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _698_
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _699_
timestamp 0
transform -1 0 9476 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _700_
timestamp 0
transform 1 0 7360 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _701_
timestamp 0
transform 1 0 7820 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _702_
timestamp 0
transform 1 0 8280 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _703_
timestamp 0
transform 1 0 6532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _704_
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _705_
timestamp 0
transform 1 0 5520 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _706_
timestamp 0
transform 1 0 6808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _707_
timestamp 0
transform -1 0 7084 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _708_
timestamp 0
transform -1 0 7452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _709_
timestamp 0
transform -1 0 9936 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _710_
timestamp 0
transform 1 0 9844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _711_
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _712_
timestamp 0
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _713_
timestamp 0
transform -1 0 8556 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _714_
timestamp 0
transform -1 0 9384 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _715_
timestamp 0
transform -1 0 8096 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _716_
timestamp 0
transform 1 0 7452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _717_
timestamp 0
transform 1 0 7820 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _718_
timestamp 0
transform -1 0 7544 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _719_
timestamp 0
transform 1 0 5060 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _720_
timestamp 0
transform 1 0 7084 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _721_
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _722_
timestamp 0
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _723_
timestamp 0
transform 1 0 5336 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _724_
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_2  _725_
timestamp 0
transform 1 0 6348 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _726_
timestamp 0
transform -1 0 6256 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _727_
timestamp 0
transform -1 0 6256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _728_
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _729_
timestamp 0
transform -1 0 9476 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _730_
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _731_
timestamp 0
transform 1 0 6808 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _732_
timestamp 0
transform -1 0 7360 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _733_
timestamp 0
transform -1 0 9292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _734_
timestamp 0
transform 1 0 7912 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _735_
timestamp 0
transform 1 0 6624 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _736_
timestamp 0
transform -1 0 6992 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _737_
timestamp 0
transform -1 0 7544 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_4  _738_
timestamp 0
transform 1 0 6900 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__o22ai_1  _739_
timestamp 0
transform -1 0 7728 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _740_
timestamp 0
transform 1 0 7728 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _741_
timestamp 0
transform -1 0 8740 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _742_
timestamp 0
transform -1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _743_
timestamp 0
transform 1 0 7728 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _744_
timestamp 0
transform 1 0 7084 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _745_
timestamp 0
transform -1 0 5612 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _746_
timestamp 0
transform 1 0 5704 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _747_
timestamp 0
transform 1 0 5980 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _748_
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a311oi_1  _749_
timestamp 0
transform -1 0 6256 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _750_
timestamp 0
transform -1 0 11960 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _751_
timestamp 0
transform -1 0 10948 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _752_
timestamp 0
transform 1 0 3956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _753_
timestamp 0
transform -1 0 8096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _754_
timestamp 0
transform 1 0 5244 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _755_
timestamp 0
transform 1 0 5336 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _756_
timestamp 0
transform -1 0 6164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _757_
timestamp 0
transform -1 0 4324 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _758_
timestamp 0
transform -1 0 5336 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _759_
timestamp 0
transform -1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _760_
timestamp 0
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _761_
timestamp 0
transform -1 0 6716 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _762_
timestamp 0
transform 1 0 5060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _763_
timestamp 0
transform 1 0 4508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _764_
timestamp 0
transform -1 0 5796 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _765_
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _766_
timestamp 0
transform 1 0 4416 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _767_
timestamp 0
transform -1 0 6808 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _768_
timestamp 0
transform -1 0 6164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _769_
timestamp 0
transform 1 0 4968 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _770_
timestamp 0
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _771_
timestamp 0
transform -1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _772_
timestamp 0
transform 1 0 16100 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _773_
timestamp 0
transform -1 0 16560 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _774_
timestamp 0
transform -1 0 17388 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _775_
timestamp 0
transform -1 0 16928 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _776_
timestamp 0
transform -1 0 16192 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _777_
timestamp 0
transform -1 0 15456 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _778_
timestamp 0
transform 1 0 13340 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _779_
timestamp 0
transform 1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _780_
timestamp 0
transform 1 0 12144 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _781_
timestamp 0
transform 1 0 12328 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _782_
timestamp 0
transform -1 0 11960 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _783_
timestamp 0
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _784_
timestamp 0
transform 1 0 9568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _785_
timestamp 0
transform -1 0 11040 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _786_
timestamp 0
transform 1 0 10120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _787_
timestamp 0
transform -1 0 15548 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _788_
timestamp 0
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _789_
timestamp 0
transform 1 0 7084 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _790_
timestamp 0
transform -1 0 7820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _791_
timestamp 0
transform 1 0 5520 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _792_
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _793_
timestamp 0
transform -1 0 5428 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _794_
timestamp 0
transform 1 0 5060 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _795_
timestamp 0
transform 1 0 3496 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _796_
timestamp 0
transform 1 0 4508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _797_
timestamp 0
transform -1 0 3128 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _798_
timestamp 0
transform -1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _799_
timestamp 0
transform -1 0 2668 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _800_
timestamp 0
transform 1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _801_
timestamp 0
transform -1 0 2576 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _802_
timestamp 0
transform -1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _803_
timestamp 0
transform 1 0 1748 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _804_
timestamp 0
transform 1 0 2208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _805_
timestamp 0
transform 1 0 9844 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _806_
timestamp 0
transform 1 0 10304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _807_
timestamp 0
transform 1 0 15456 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _808_
timestamp 0
transform 1 0 15272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _809_
timestamp 0
transform -1 0 15272 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _810_
timestamp 0
transform -1 0 16468 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _811_
timestamp 0
transform -1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _812_
timestamp 0
transform 1 0 15824 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _813_
timestamp 0
transform 1 0 14904 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _814_
timestamp 0
transform 1 0 14904 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _815_
timestamp 0
transform 1 0 15364 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _816_
timestamp 0
transform -1 0 15824 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _817_
timestamp 0
transform -1 0 13708 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _818_
timestamp 0
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _819_
timestamp 0
transform -1 0 13248 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _820_
timestamp 0
transform -1 0 12420 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _821_
timestamp 0
transform -1 0 15180 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _822_
timestamp 0
transform 1 0 15180 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _823_
timestamp 0
transform -1 0 14904 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _824_
timestamp 0
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _825_
timestamp 0
transform 1 0 12604 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _826_
timestamp 0
transform -1 0 14812 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _827_
timestamp 0
transform -1 0 15824 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _828_
timestamp 0
transform -1 0 15640 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _829_
timestamp 0
transform -1 0 15364 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _830_
timestamp 0
transform 1 0 14444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _831_
timestamp 0
transform 1 0 14812 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _832_
timestamp 0
transform -1 0 14444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _833_
timestamp 0
transform 1 0 13708 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _834_
timestamp 0
transform -1 0 15180 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _835_
timestamp 0
transform -1 0 15272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _836_
timestamp 0
transform 1 0 14352 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _837_
timestamp 0
transform 1 0 15180 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _838_
timestamp 0
transform -1 0 15640 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _839_
timestamp 0
transform 1 0 14444 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _840_
timestamp 0
transform 1 0 16008 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _841_
timestamp 0
transform -1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _842_
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _843_
timestamp 0
transform 1 0 17388 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _844_
timestamp 0
transform 1 0 16100 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _845_
timestamp 0
transform -1 0 17664 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _846_
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _847_
timestamp 0
transform 1 0 17940 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _848_
timestamp 0
transform -1 0 17940 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _849_
timestamp 0
transform 1 0 16652 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _850_
timestamp 0
transform -1 0 16100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _851_
timestamp 0
transform -1 0 16928 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _852_
timestamp 0
transform 1 0 16376 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _853_
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _854_
timestamp 0
transform -1 0 15456 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _855_
timestamp 0
transform -1 0 16560 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _856_
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _857_
timestamp 0
transform -1 0 17664 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _858_
timestamp 0
transform -1 0 17020 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _859_
timestamp 0
transform 1 0 14996 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _860_
timestamp 0
transform 1 0 15824 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _861_
timestamp 0
transform 1 0 14352 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _862_
timestamp 0
transform -1 0 15364 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _863_
timestamp 0
transform 1 0 15364 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _864_
timestamp 0
transform -1 0 14352 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _865_
timestamp 0
transform 1 0 10856 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _866_
timestamp 0
transform -1 0 12052 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _867_
timestamp 0
transform 1 0 3128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _868_
timestamp 0
transform 1 0 5152 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _869_
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _870_
timestamp 0
transform 1 0 3128 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _871_
timestamp 0
transform 1 0 4784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _872_
timestamp 0
transform 1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _873_
timestamp 0
transform -1 0 3864 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _874_
timestamp 0
transform -1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _875_
timestamp 0
transform 1 0 2300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _876_
timestamp 0
transform -1 0 3680 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _877_
timestamp 0
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _878_
timestamp 0
transform 1 0 2852 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _879_
timestamp 0
transform -1 0 5244 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _880_
timestamp 0
transform -1 0 3128 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _881_
timestamp 0
transform 1 0 2760 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _882_
timestamp 0
transform -1 0 3864 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _883_
timestamp 0
transform -1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _884_
timestamp 0
transform 1 0 2852 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _885_
timestamp 0
transform -1 0 3588 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _886_
timestamp 0
transform 1 0 2944 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _887_
timestamp 0
transform 1 0 9016 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _888_
timestamp 0
transform -1 0 11408 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _889_
timestamp 0
transform 1 0 9844 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _890_
timestamp 0
transform 1 0 10488 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _891_
timestamp 0
transform 1 0 9660 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _892_
timestamp 0
transform 1 0 9752 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _893_
timestamp 0
transform 1 0 9936 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _894_
timestamp 0
transform 1 0 11684 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _895_
timestamp 0
transform -1 0 16376 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _896_
timestamp 0
transform 1 0 18492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _897_
timestamp 0
transform 1 0 14628 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _898_
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _899_
timestamp 0
transform 1 0 12880 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _900_
timestamp 0
transform -1 0 18124 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _901_
timestamp 0
transform -1 0 19596 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _902_
timestamp 0
transform 1 0 17020 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _903_
timestamp 0
transform -1 0 19504 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _904_
timestamp 0
transform -1 0 20976 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _905_
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _906_
timestamp 0
transform -1 0 20608 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _907_
timestamp 0
transform 1 0 20516 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _908_
timestamp 0
transform 1 0 19504 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _909_
timestamp 0
transform 1 0 18032 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _910_
timestamp 0
transform 1 0 17572 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _911_
timestamp 0
transform 1 0 20056 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _912_
timestamp 0
transform 1 0 19964 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _913_
timestamp 0
transform 1 0 10488 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _914_
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _915_
timestamp 0
transform -1 0 9844 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _916_
timestamp 0
transform -1 0 8188 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _917_
timestamp 0
transform -1 0 8372 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _918_
timestamp 0
transform 1 0 9936 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _919_
timestamp 0
transform -1 0 13248 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _920_
timestamp 0
transform 1 0 8924 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _921_
timestamp 0
transform -1 0 15364 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _922_
timestamp 0
transform -1 0 17112 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _923_
timestamp 0
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _924_
timestamp 0
transform 1 0 20516 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _925_
timestamp 0
transform -1 0 21712 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _926_
timestamp 0
transform 1 0 19596 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _927_
timestamp 0
transform 1 0 18124 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _928_
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _929_
timestamp 0
transform 1 0 16284 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _930_
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _931_
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _932_
timestamp 0
transform 1 0 13616 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _933_
timestamp 0
transform 1 0 20516 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _934_
timestamp 0
transform 1 0 20240 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _935_
timestamp 0
transform 1 0 19872 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _936_
timestamp 0
transform 1 0 18400 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _937_
timestamp 0
transform 1 0 16928 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _938_
timestamp 0
transform -1 0 18124 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _939_
timestamp 0
transform 1 0 17020 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _940_
timestamp 0
transform -1 0 20700 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _941_
timestamp 0
transform 1 0 13984 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _942_
timestamp 0
transform 1 0 5336 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _943_
timestamp 0
transform 1 0 7084 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _944_
timestamp 0
transform 1 0 7176 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _945_
timestamp 0
transform 1 0 4600 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _946_
timestamp 0
transform 1 0 4876 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _947_
timestamp 0
transform 1 0 7360 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _948_
timestamp 0
transform -1 0 9476 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _949_
timestamp 0
transform 1 0 5152 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _950_
timestamp 0
transform -1 0 11408 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _951_
timestamp 0
transform 1 0 3128 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _952_
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _953_
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _954_
timestamp 0
transform -1 0 5612 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _955_
timestamp 0
transform 1 0 4048 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _956_
timestamp 0
transform 1 0 4416 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _957_
timestamp 0
transform 1 0 4968 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _958_
timestamp 0
transform -1 0 8280 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _959_
timestamp 0
transform 1 0 7636 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _960_
timestamp 0
transform -1 0 17480 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _961_
timestamp 0
transform -1 0 18400 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _962_
timestamp 0
transform 1 0 15456 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _963_
timestamp 0
transform 1 0 13800 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _964_
timestamp 0
transform 1 0 11868 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _965_
timestamp 0
transform 1 0 10396 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _966_
timestamp 0
transform 1 0 9936 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _967_
timestamp 0
transform -1 0 15548 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _968_
timestamp 0
transform 1 0 20424 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _969_
timestamp 0
transform -1 0 8556 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _970_
timestamp 0
transform 1 0 4784 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _971_
timestamp 0
transform 1 0 4600 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _972_
timestamp 0
transform 1 0 4048 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _973_
timestamp 0
transform 1 0 2024 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _974_
timestamp 0
transform 1 0 1472 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _975_
timestamp 0
transform 1 0 2116 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _976_
timestamp 0
transform 1 0 1564 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _977_
timestamp 0
transform 1 0 9108 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _978_
timestamp 0
transform 1 0 12420 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _979_
timestamp 0
transform 1 0 12052 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _980_
timestamp 0
transform 1 0 14812 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _981_
timestamp 0
transform -1 0 13984 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _982_
timestamp 0
transform 1 0 16284 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _983_
timestamp 0
transform -1 0 19136 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _984_
timestamp 0
transform -1 0 17940 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _985_
timestamp 0
transform -1 0 15548 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _986_
timestamp 0
transform 1 0 12144 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _987_
timestamp 0
transform 1 0 3404 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _988_
timestamp 0
transform 1 0 2024 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _989_
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _990_
timestamp 0
transform 1 0 1656 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _991_
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _992_
timestamp 0
transform 1 0 2208 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _993_
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _994_
timestamp 0
transform 1 0 2668 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 11684 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 0
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 0
transform 1 0 5244 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 0
transform -1 0 4416 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 0
transform -1 0 9660 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 0
transform -1 0 14812 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 0
transform 1 0 18216 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 0
transform 1 0 15640 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 0
transform 1 0 18216 0 -1 13056
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6
timestamp 0
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18
timestamp 0
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26
timestamp 0
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_91
timestamp 0
transform 1 0 9476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_103
timestamp 0
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 0
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_136
timestamp 0
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_175
timestamp 0
transform 1 0 17204 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_182
timestamp 0
transform 1 0 17848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_194
timestamp 0
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_200
timestamp 0
transform 1 0 19504 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_212
timestamp 0
transform 1 0 20608 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_220
timestamp 0
transform 1 0 21344 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_35
timestamp 0
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_82
timestamp 0
transform 1 0 8648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_104
timestamp 0
transform 1 0 10672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_124
timestamp 0
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_144
timestamp 0
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 0
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_201
timestamp 0
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_210
timestamp 0
transform 1 0 20424 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_222
timestamp 0
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_225
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_58
timestamp 0
transform 1 0 6440 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_72
timestamp 0
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_99
timestamp 0
transform 1 0 10212 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_171
timestamp 0
transform 1 0 16836 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_208
timestamp 0
transform 1 0 20240 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_220
timestamp 0
transform 1 0 21344 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_226
timestamp 0
transform 1 0 21896 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_35
timestamp 0
transform 1 0 4324 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_65
timestamp 0
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_80
timestamp 0
transform 1 0 8464 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_88
timestamp 0
transform 1 0 9200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_99
timestamp 0
transform 1 0 10212 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_135
timestamp 0
transform 1 0 13524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_151
timestamp 0
transform 1 0 14996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 0
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_174
timestamp 0
transform 1 0 17112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_216
timestamp 0
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_225
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_45
timestamp 0
transform 1 0 5244 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_51
timestamp 0
transform 1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_56
timestamp 0
transform 1 0 6256 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_64
timestamp 0
transform 1 0 6992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_76
timestamp 0
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_121
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_129
timestamp 0
transform 1 0 12972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_154
timestamp 0
transform 1 0 15272 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_167
timestamp 0
transform 1 0 16468 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_192
timestamp 0
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 0
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 0
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_221
timestamp 0
transform 1 0 21436 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_35
timestamp 0
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_46
timestamp 0
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 0
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_63
timestamp 0
transform 1 0 6900 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_74
timestamp 0
transform 1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_80
timestamp 0
transform 1 0 8464 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_92
timestamp 0
transform 1 0 9568 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_97
timestamp 0
transform 1 0 10028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 0
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_149
timestamp 0
transform 1 0 14812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_153
timestamp 0
transform 1 0 15180 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166
timestamp 0
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_177
timestamp 0
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_184
timestamp 0
transform 1 0 18032 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_216
timestamp 0
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_225
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_61
timestamp 0
transform 1 0 6716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_79
timestamp 0
transform 1 0 8372 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_89
timestamp 0
transform 1 0 9292 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_122
timestamp 0
transform 1 0 12328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_129
timestamp 0
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 0
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_157
timestamp 0
transform 1 0 15548 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_168
timestamp 0
transform 1 0 16560 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_180
timestamp 0
transform 1 0 17664 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_192
timestamp 0
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_197
timestamp 0
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_211
timestamp 0
transform 1 0 20516 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_220
timestamp 0
transform 1 0 21344 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_226
timestamp 0
transform 1 0 21896 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_52
timestamp 0
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_68
timestamp 0
transform 1 0 7360 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_83
timestamp 0
transform 1 0 8740 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_123
timestamp 0
transform 1 0 12420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_137
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_158
timestamp 0
transform 1 0 15640 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 0
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 0
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_225
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_46
timestamp 0
transform 1 0 5336 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_58
timestamp 0
transform 1 0 6440 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_70
timestamp 0
transform 1 0 7544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_74
timestamp 0
transform 1 0 7912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_79
timestamp 0
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_106
timestamp 0
transform 1 0 10856 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_119
timestamp 0
transform 1 0 12052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_131
timestamp 0
transform 1 0 13156 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_150
timestamp 0
transform 1 0 14904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_157
timestamp 0
transform 1 0 15548 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 0
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_207
timestamp 0
transform 1 0 20148 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_36
timestamp 0
transform 1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_44
timestamp 0
transform 1 0 5152 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 0
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_72
timestamp 0
transform 1 0 7728 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_77
timestamp 0
transform 1 0 8188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_89
timestamp 0
transform 1 0 9292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_101
timestamp 0
transform 1 0 10396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_109
timestamp 0
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_120
timestamp 0
transform 1 0 12144 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_132
timestamp 0
transform 1 0 13248 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_150
timestamp 0
transform 1 0 14904 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_162
timestamp 0
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_179
timestamp 0
transform 1 0 17572 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_207
timestamp 0
transform 1 0 20148 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_225
timestamp 0
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_76
timestamp 0
transform 1 0 8096 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 0
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_93
timestamp 0
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_99
timestamp 0
transform 1 0 10212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_118
timestamp 0
transform 1 0 11960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_128
timestamp 0
transform 1 0 12880 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_136
timestamp 0
transform 1 0 13616 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_149
timestamp 0
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_157
timestamp 0
transform 1 0 15548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_161
timestamp 0
transform 1 0 15916 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_181
timestamp 0
transform 1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_192
timestamp 0
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_200
timestamp 0
transform 1 0 19504 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_206
timestamp 0
transform 1 0 20056 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_226
timestamp 0
transform 1 0 21896 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_21
timestamp 0
transform 1 0 3036 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_38
timestamp 0
transform 1 0 4600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_65
timestamp 0
transform 1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_129
timestamp 0
transform 1 0 12972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_133
timestamp 0
transform 1 0 13340 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_156
timestamp 0
transform 1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_164
timestamp 0
transform 1 0 16192 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 0
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_205
timestamp 0
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_213
timestamp 0
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 0
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_225
timestamp 0
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_6
timestamp 0
transform 1 0 1656 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_43
timestamp 0
transform 1 0 5060 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_60
timestamp 0
transform 1 0 6624 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_128
timestamp 0
transform 1 0 12880 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_157
timestamp 0
transform 1 0 15548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_169
timestamp 0
transform 1 0 16652 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_178
timestamp 0
transform 1 0 17480 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_190
timestamp 0
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_21
timestamp 0
transform 1 0 3036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_29
timestamp 0
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_34
timestamp 0
transform 1 0 4232 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_42
timestamp 0
transform 1 0 4968 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_68
timestamp 0
transform 1 0 7360 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_74
timestamp 0
transform 1 0 7912 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_102
timestamp 0
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 0
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_117
timestamp 0
transform 1 0 11868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_129
timestamp 0
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_138
timestamp 0
transform 1 0 13800 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_150
timestamp 0
transform 1 0 14904 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_162
timestamp 0
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_177
timestamp 0
transform 1 0 17388 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_185
timestamp 0
transform 1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_220
timestamp 0
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_225
timestamp 0
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_7
timestamp 0
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_55
timestamp 0
transform 1 0 6164 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_62
timestamp 0
transform 1 0 6808 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_74
timestamp 0
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 0
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_91
timestamp 0
transform 1 0 9476 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_103
timestamp 0
transform 1 0 10580 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_115
timestamp 0
transform 1 0 11684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_119
timestamp 0
transform 1 0 12052 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_125
timestamp 0
transform 1 0 12604 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_129
timestamp 0
transform 1 0 12972 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_136
timestamp 0
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_152
timestamp 0
transform 1 0 15088 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_172
timestamp 0
transform 1 0 16928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_182
timestamp 0
transform 1 0 17848 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_224
timestamp 0
transform 1 0 21712 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_32
timestamp 0
transform 1 0 4048 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_76
timestamp 0
transform 1 0 8096 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_88
timestamp 0
transform 1 0 9200 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_118
timestamp 0
transform 1 0 11960 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_135
timestamp 0
transform 1 0 13524 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_164
timestamp 0
transform 1 0 16192 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_188
timestamp 0
transform 1 0 18400 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_225
timestamp 0
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_36
timestamp 0
transform 1 0 4416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_54
timestamp 0
transform 1 0 6072 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 0
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_91
timestamp 0
transform 1 0 9476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_96
timestamp 0
transform 1 0 9936 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_178
timestamp 0
transform 1 0 17480 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_190
timestamp 0
transform 1 0 18584 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_215
timestamp 0
transform 1 0 20884 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_20
timestamp 0
transform 1 0 2944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_30
timestamp 0
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_62
timestamp 0
transform 1 0 6808 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_83
timestamp 0
transform 1 0 8740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_108
timestamp 0
transform 1 0 11040 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_177
timestamp 0
transform 1 0 17388 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_183
timestamp 0
transform 1 0 17940 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_208
timestamp 0
transform 1 0 20240 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_220
timestamp 0
transform 1 0 21344 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_225
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_9
timestamp 0
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 0
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_40
timestamp 0
transform 1 0 4784 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_46
timestamp 0
transform 1 0 5336 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_56
timestamp 0
transform 1 0 6256 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_68
timestamp 0
transform 1 0 7360 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_80
timestamp 0
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_103
timestamp 0
transform 1 0 10580 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_111
timestamp 0
transform 1 0 11316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_115
timestamp 0
transform 1 0 11684 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_119
timestamp 0
transform 1 0 12052 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_131
timestamp 0
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_146
timestamp 0
transform 1 0 14536 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_158
timestamp 0
transform 1 0 15640 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_170
timestamp 0
transform 1 0 16744 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 0
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_222
timestamp 0
transform 1 0 21528 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_226
timestamp 0
transform 1 0 21896 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_23
timestamp 0
transform 1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_31
timestamp 0
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_43
timestamp 0
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_61
timestamp 0
transform 1 0 6716 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_135
timestamp 0
transform 1 0 13524 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_147
timestamp 0
transform 1 0 14628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_159
timestamp 0
transform 1 0 15732 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_222
timestamp 0
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_225
timestamp 0
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_45
timestamp 0
transform 1 0 5244 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_62
timestamp 0
transform 1 0 6808 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_67
timestamp 0
transform 1 0 7268 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 0
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_91
timestamp 0
transform 1 0 9476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_111
timestamp 0
transform 1 0 11316 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_119
timestamp 0
transform 1 0 12052 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_136
timestamp 0
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_157
timestamp 0
transform 1 0 15548 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_174
timestamp 0
transform 1 0 17112 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_186
timestamp 0
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 0
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_224
timestamp 0
transform 1 0 21712 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_15
timestamp 0
transform 1 0 2484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_21
timestamp 0
transform 1 0 3036 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_41
timestamp 0
transform 1 0 4876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_118
timestamp 0
transform 1 0 11960 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_135
timestamp 0
transform 1 0 13524 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_143
timestamp 0
transform 1 0 14260 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_173
timestamp 0
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_190
timestamp 0
transform 1 0 18584 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_202
timestamp 0
transform 1 0 19688 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_221
timestamp 0
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 0
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_9
timestamp 0
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 0
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_57
timestamp 0
transform 1 0 6348 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_98
timestamp 0
transform 1 0 10120 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_107
timestamp 0
transform 1 0 10948 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_113
timestamp 0
transform 1 0 11500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_135
timestamp 0
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_145
timestamp 0
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_160
timestamp 0
transform 1 0 15824 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 0
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 0
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 0
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_221
timestamp 0
transform 1 0 21436 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_19
timestamp 0
transform 1 0 2852 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_44
timestamp 0
transform 1 0 5152 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_63
timestamp 0
transform 1 0 6900 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_75
timestamp 0
transform 1 0 8004 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_87
timestamp 0
transform 1 0 9108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_99
timestamp 0
transform 1 0 10212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_119
timestamp 0
transform 1 0 12052 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_139
timestamp 0
transform 1 0 13892 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_149
timestamp 0
transform 1 0 14812 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_159
timestamp 0
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_185
timestamp 0
transform 1 0 18124 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_216
timestamp 0
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_225
timestamp 0
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_11
timestamp 0
transform 1 0 2116 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_46
timestamp 0
transform 1 0 5336 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_58
timestamp 0
transform 1 0 6440 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_66
timestamp 0
transform 1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_80
timestamp 0
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 0
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_121
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_156
timestamp 0
transform 1 0 15456 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_202
timestamp 0
transform 1 0 19688 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_209
timestamp 0
transform 1 0 20332 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_11
timestamp 0
transform 1 0 2116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_62
timestamp 0
transform 1 0 6808 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_93
timestamp 0
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_131
timestamp 0
transform 1 0 13156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_139
timestamp 0
transform 1 0 13892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_165
timestamp 0
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_196
timestamp 0
transform 1 0 19136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_203
timestamp 0
transform 1 0 19780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_225
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_22
timestamp 0
transform 1 0 3128 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_37
timestamp 0
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_54
timestamp 0
transform 1 0 6072 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 0
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_90
timestamp 0
transform 1 0 9384 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_119
timestamp 0
transform 1 0 12052 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_135
timestamp 0
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_160
timestamp 0
transform 1 0 15824 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_172
timestamp 0
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_176
timestamp 0
transform 1 0 17296 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_197
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_224
timestamp 0
transform 1 0 21712 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_39
timestamp 0
transform 1 0 4692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_50
timestamp 0
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_61
timestamp 0
transform 1 0 6716 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_81
timestamp 0
transform 1 0 8556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_85
timestamp 0
transform 1 0 8924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_102
timestamp 0
transform 1 0 10488 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_121
timestamp 0
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_135
timestamp 0
transform 1 0 13524 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_143
timestamp 0
transform 1 0 14260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_158
timestamp 0
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 0
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_187
timestamp 0
transform 1 0 18308 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_220
timestamp 0
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_225
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_15
timestamp 0
transform 1 0 2484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_23
timestamp 0
transform 1 0 3220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_37
timestamp 0
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_43
timestamp 0
transform 1 0 5060 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_55
timestamp 0
transform 1 0 6164 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_67
timestamp 0
transform 1 0 7268 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_79
timestamp 0
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_93
timestamp 0
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_121
timestamp 0
transform 1 0 12236 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_130
timestamp 0
transform 1 0 13064 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 0
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_158
timestamp 0
transform 1 0 15640 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_181
timestamp 0
transform 1 0 17756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_193
timestamp 0
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 0
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_201
timestamp 0
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_205
timestamp 0
transform 1 0 19964 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_213
timestamp 0
transform 1 0 20700 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_223
timestamp 0
transform 1 0 21620 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_15
timestamp 0
transform 1 0 2484 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_24
timestamp 0
transform 1 0 3312 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_45
timestamp 0
transform 1 0 5244 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_91
timestamp 0
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_133
timestamp 0
transform 1 0 13340 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_154
timestamp 0
transform 1 0 15272 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 0
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_179
timestamp 0
transform 1 0 17572 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_191
timestamp 0
transform 1 0 18676 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_203
timestamp 0
transform 1 0 19780 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_215
timestamp 0
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 0
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_11
timestamp 0
transform 1 0 2116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_57
timestamp 0
transform 1 0 6348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_89
timestamp 0
transform 1 0 9292 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_95
timestamp 0
transform 1 0 9844 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_123
timestamp 0
transform 1 0 12420 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_164
timestamp 0
transform 1 0 16192 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_168
timestamp 0
transform 1 0 16560 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_172
timestamp 0
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_176
timestamp 0
transform 1 0 17296 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_187
timestamp 0
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 0
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_213
timestamp 0
transform 1 0 20700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_225
timestamp 0
transform 1 0 21804 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_30
timestamp 0
transform 1 0 3864 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_42
timestamp 0
transform 1 0 4968 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_50
timestamp 0
transform 1 0 5704 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_70
timestamp 0
transform 1 0 7544 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_80
timestamp 0
transform 1 0 8464 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_92
timestamp 0
transform 1 0 9568 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_103
timestamp 0
transform 1 0 10580 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 0
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_113
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_135
timestamp 0
transform 1 0 13524 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_147
timestamp 0
transform 1 0 14628 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_159
timestamp 0
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_199
timestamp 0
transform 1 0 19412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_211
timestamp 0
transform 1 0 20516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 0
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_225
timestamp 0
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_15
timestamp 0
transform 1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_25
timestamp 0
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_43
timestamp 0
transform 1 0 5060 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_55
timestamp 0
transform 1 0 6164 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_67
timestamp 0
transform 1 0 7268 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_79
timestamp 0
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 0
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 0
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 0
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_121
timestamp 0
transform 1 0 12236 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 0
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_153
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_160
timestamp 0
transform 1 0 15824 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_172
timestamp 0
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_176
timestamp 0
transform 1 0 17296 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_184
timestamp 0
transform 1 0 18032 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_202
timestamp 0
transform 1 0 19688 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_211
timestamp 0
transform 1 0 20516 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_223
timestamp 0
transform 1 0 21620 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_15
timestamp 0
transform 1 0 2484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_23
timestamp 0
transform 1 0 3220 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_31
timestamp 0
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_43
timestamp 0
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 0
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_64
timestamp 0
transform 1 0 6992 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_76
timestamp 0
transform 1 0 8096 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_84
timestamp 0
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_91
timestamp 0
transform 1 0 9476 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_110
timestamp 0
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_117
timestamp 0
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_122
timestamp 0
transform 1 0 12328 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_126
timestamp 0
transform 1 0 12696 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_138
timestamp 0
transform 1 0 13800 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_150
timestamp 0
transform 1 0 14904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 0
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_173
timestamp 0
transform 1 0 17020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_185
timestamp 0
transform 1 0 18124 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_197
timestamp 0
transform 1 0 19228 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_205
timestamp 0
transform 1 0 19964 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_212
timestamp 0
transform 1 0 20608 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_225
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 0
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_15
timestamp 0
transform 1 0 2484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 0
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_36
timestamp 0
transform 1 0 4416 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_48
timestamp 0
transform 1 0 5520 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_58
timestamp 0
transform 1 0 6440 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 0
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_85
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_123
timestamp 0
transform 1 0 12420 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_135
timestamp 0
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 0
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_147
timestamp 0
transform 1 0 14628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_162
timestamp 0
transform 1 0 16008 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_168
timestamp 0
transform 1 0 16560 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_174
timestamp 0
transform 1 0 17112 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_186
timestamp 0
transform 1 0 18216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 0
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 0
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_221
timestamp 0
transform 1 0 21436 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_3
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_11
timestamp 0
transform 1 0 2116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_33
timestamp 0
transform 1 0 4140 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_41
timestamp 0
transform 1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_73
timestamp 0
transform 1 0 7820 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_91
timestamp 0
transform 1 0 9476 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_99
timestamp 0
transform 1 0 10212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_110
timestamp 0
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_156
timestamp 0
transform 1 0 15456 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_180
timestamp 0
transform 1 0 17664 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_192
timestamp 0
transform 1 0 18768 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_204
timestamp 0
transform 1 0 19872 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_216
timestamp 0
transform 1 0 20976 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_220
timestamp 0
transform 1 0 21344 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_225
timestamp 0
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_15
timestamp 0
transform 1 0 2484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_19
timestamp 0
transform 1 0 2852 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_24
timestamp 0
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_37
timestamp 0
transform 1 0 4508 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_43
timestamp 0
transform 1 0 5060 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_60
timestamp 0
transform 1 0 6624 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_66
timestamp 0
transform 1 0 7176 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_75
timestamp 0
transform 1 0 8004 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 0
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_93
timestamp 0
transform 1 0 9660 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 0
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_157
timestamp 0
transform 1 0 15548 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_165
timestamp 0
transform 1 0 16284 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_183
timestamp 0
transform 1 0 17940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 0
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 0
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_221
timestamp 0
transform 1 0 21436 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_9
timestamp 0
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_21
timestamp 0
transform 1 0 3036 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_27
timestamp 0
transform 1 0 3588 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_29
timestamp 0
transform 1 0 3772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_41
timestamp 0
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_53
timestamp 0
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 0
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_81
timestamp 0
transform 1 0 8556 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_85
timestamp 0
transform 1 0 8924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_97
timestamp 0
transform 1 0 10028 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_107
timestamp 0
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 0
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_125
timestamp 0
transform 1 0 12604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_131
timestamp 0
transform 1 0 13156 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_138
timestamp 0
transform 1 0 13800 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_141
timestamp 0
transform 1 0 14076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_153
timestamp 0
transform 1 0 15180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_165
timestamp 0
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_169
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_173
timestamp 0
transform 1 0 17020 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_185
timestamp 0
transform 1 0 18124 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_193
timestamp 0
transform 1 0 18860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_197
timestamp 0
transform 1 0 19228 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_202
timestamp 0
transform 1 0 19688 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_214
timestamp 0
transform 1 0 20792 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 0
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 4508 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform 1 0 7360 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform -1 0 5336 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 11868 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform -1 0 4508 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform -1 0 5060 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform -1 0 12144 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform -1 0 12236 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform -1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform -1 0 6256 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform -1 0 17572 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 0
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 0
transform -1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 0
transform -1 0 11408 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 0
transform -1 0 11132 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 0
transform -1 0 11960 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 0
transform -1 0 4140 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 0
transform -1 0 12052 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 0
transform -1 0 12328 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 0
transform -1 0 16284 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 0
transform -1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 0
transform -1 0 5888 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold27
timestamp 0
transform 1 0 6992 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 0
transform 1 0 6348 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 0
transform -1 0 6256 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold30
timestamp 0
transform -1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 0
transform -1 0 4600 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 0
transform 1 0 18032 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 0
transform 1 0 19504 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 0
transform 1 0 19504 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 0
transform -1 0 4048 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 0
transform -1 0 3864 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 0
transform -1 0 19136 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 0
transform 1 0 20424 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 0
transform -1 0 18676 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 0
transform 1 0 15272 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 0
transform -1 0 21712 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 0
transform -1 0 14812 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 0
transform -1 0 4508 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 0
transform 1 0 18400 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 0
transform -1 0 12604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 0
transform -1 0 18768 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 0
transform -1 0 21620 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 0
transform -1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 0
transform -1 0 6256 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 0
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 0
transform -1 0 21620 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 0
transform -1 0 6624 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 0
transform -1 0 21712 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 0
transform -1 0 19964 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 0
transform -1 0 3312 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 0
transform -1 0 12788 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 0
transform 1 0 17480 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 0
transform -1 0 20516 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 0
transform -1 0 19964 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 0
transform -1 0 20516 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 0
transform -1 0 18860 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 0
transform -1 0 14996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 0
transform -1 0 21344 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 0
transform -1 0 18676 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 0
transform -1 0 13524 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 0
transform -1 0 4508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 0
transform -1 0 15916 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 0
transform -1 0 17848 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 0
transform -1 0 18584 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 0
transform -1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 0
transform -1 0 14812 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 0
transform -1 0 6164 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 0
transform -1 0 11776 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 0
transform -1 0 7820 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 0
transform -1 0 18676 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 0
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 0
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform 1 0 19412 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 0
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 0
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform -1 0 21712 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 0
transform -1 0 1932 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform -1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 22264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 22264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 22264 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 22264 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 22264 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 22264 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 22264 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 22264 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 22264 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 22264 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 22264 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 22264 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 22264 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 22264 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 22264 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 22264 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 22264 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 22264 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 22264 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 0
transform -1 0 22264 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 0
transform -1 0 22264 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 0
transform -1 0 22264 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 0
transform -1 0 22264 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 0
transform -1 0 22264 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 0
transform -1 0 22264 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 0
transform -1 0 22264 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 0
transform -1 0 22264 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 0
transform -1 0 22264 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 0
transform -1 0 22264 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 0
transform -1 0 22264 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 0
transform 1 0 3680 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 0
transform 1 0 8832 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 0
transform 1 0 13984 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 0
transform 1 0 19136 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
<< labels >>
rlabel metal1 s 11684 22848 11684 22848 4 VGND
rlabel metal1 s 11684 22304 11684 22304 4 VPWR
rlabel metal1 s 16146 4726 16146 4726 4 _000_
rlabel metal1 s 16238 4794 16238 4794 4 _001_
rlabel metal1 s 19044 7378 19044 7378 4 _002_
rlabel metal1 s 18492 7310 18492 7310 4 _003_
rlabel metal1 s 19550 14926 19550 14926 4 _004_
rlabel metal1 s 19274 14484 19274 14484 4 _005_
rlabel metal1 s 13938 11764 13938 11764 4 _006_
rlabel metal1 s 13616 11662 13616 11662 4 _007_
rlabel metal1 s 8004 11730 8004 11730 4 _008_
rlabel metal1 s 7636 11662 7636 11662 4 _009_
rlabel metal1 s 20792 11730 20792 11730 4 _010_
rlabel metal2 s 21022 11968 21022 11968 4 _011_
rlabel metal2 s 9323 17170 9323 17170 4 _012_
rlabel metal1 s 12512 15946 12512 15946 4 _013_
rlabel metal1 s 9966 16490 9966 16490 4 _014_
rlabel metal2 s 11270 18530 11270 18530 4 _015_
rlabel metal1 s 10115 18258 10115 18258 4 _016_
rlabel metal2 s 10258 20706 10258 20706 4 _017_
rlabel metal2 s 10442 21794 10442 21794 4 _018_
rlabel metal1 s 12047 21590 12047 21590 4 _019_
rlabel metal1 s 15543 3094 15543 3094 4 _020_
rlabel metal1 s 13922 3434 13922 3434 4 _021_
rlabel metal1 s 13294 2618 13294 2618 4 _022_
rlabel metal1 s 17342 2618 17342 2618 4 _023_
rlabel metal1 s 19094 3026 19094 3026 4 _024_
rlabel metal1 s 17142 4522 17142 4522 4 _025_
rlabel metal1 s 18956 4182 18956 4182 4 _026_
rlabel metal2 s 20194 3910 20194 3910 4 _027_
rlabel metal1 s 19228 9418 19228 9418 4 _028_
rlabel metal2 s 20470 9350 20470 9350 4 _029_
rlabel metal1 s 20971 8942 20971 8942 4 _030_
rlabel metal1 s 19580 10710 19580 10710 4 _031_
rlabel metal1 s 18809 11798 18809 11798 4 _032_
rlabel metal1 s 17694 12138 17694 12138 4 _033_
rlabel metal1 s 20276 12818 20276 12818 4 _034_
rlabel metal2 s 20281 13906 20281 13906 4 _035_
rlabel metal1 s 10518 7786 10518 7786 4 _036_
rlabel metal1 s 11720 8466 11720 8466 4 _037_
rlabel metal1 s 9434 9622 9434 9622 4 _038_
rlabel metal1 s 8065 8874 8065 8874 4 _039_
rlabel metal2 s 8065 5610 8065 5610 4 _040_
rlabel metal1 s 10345 6358 10345 6358 4 _041_
rlabel metal1 s 12332 4114 12332 4114 4 _042_
rlabel metal1 s 9655 3094 9655 3094 4 _043_
rlabel metal1 s 15241 6358 15241 6358 4 _044_
rlabel metal2 s 16514 13090 16514 13090 4 _045_
rlabel metal2 s 20833 6766 20833 6766 4 _046_
rlabel metal1 s 21492 7378 21492 7378 4 _047_
rlabel metal2 s 20286 6086 20286 6086 4 _048_
rlabel metal1 s 18625 6290 18625 6290 4 _049_
rlabel metal1 s 16866 8534 16866 8534 4 _050_
rlabel metal1 s 16406 7786 16406 7786 4 _051_
rlabel metal2 s 16054 6052 16054 6052 4 _052_
rlabel metal2 s 13846 5202 13846 5202 4 _053_
rlabel metal2 s 20930 15266 20930 15266 4 _054_
rlabel metal1 s 20362 16150 20362 16150 4 _055_
rlabel metal1 s 20040 17238 20040 17238 4 _056_
rlabel metal1 s 18216 16762 18216 16762 4 _057_
rlabel metal2 s 17245 16082 17245 16082 4 _058_
rlabel metal1 s 17904 14994 17904 14994 4 _059_
rlabel metal2 s 17618 14042 17618 14042 4 _060_
rlabel metal1 s 20152 18666 20152 18666 4 _061_
rlabel metal1 s 14030 8058 14030 8058 4 _062_
rlabel metal1 s 5837 13294 5837 13294 4 _063_
rlabel metal1 s 7360 12954 7360 12954 4 _064_
rlabel metal2 s 7493 16558 7493 16558 4 _065_
rlabel metal2 s 5750 16354 5750 16354 4 _066_
rlabel metal2 s 6394 18530 6394 18530 4 _067_
rlabel metal1 s 7815 18734 7815 18734 4 _068_
rlabel metal2 s 8510 21726 8510 21726 4 _069_
rlabel metal2 s 5750 21794 5750 21794 4 _070_
rlabel metal1 s 10998 13974 10998 13974 4 _071_
rlabel metal1 s 3721 8534 3721 8534 4 _072_
rlabel metal1 s 5147 8534 5147 8534 4 _073_
rlabel metal1 s 4135 7786 4135 7786 4 _074_
rlabel metal1 s 5535 6358 5535 6358 4 _075_
rlabel metal1 s 4600 5338 4600 5338 4 _076_
rlabel metal1 s 4682 3026 4682 3026 4 _077_
rlabel metal1 s 5182 3434 5182 3434 4 _078_
rlabel metal1 s 8065 3094 8065 3094 4 _079_
rlabel metal1 s 16698 10438 16698 10438 4 _080_
rlabel metal1 s 17484 10710 17484 10710 4 _081_
rlabel metal1 s 15578 9962 15578 9962 4 _082_
rlabel metal2 s 14858 10438 14858 10438 4 _083_
rlabel metal1 s 12277 11050 12277 11050 4 _084_
rlabel metal1 s 10943 11050 10943 11050 4 _085_
rlabel metal1 s 10253 10710 10253 10710 4 _086_
rlabel metal1 s 14996 8058 14996 8058 4 _087_
rlabel metal2 s 7774 10914 7774 10914 4 _088_
rlabel metal1 s 5561 10710 5561 10710 4 _089_
rlabel metal2 s 4917 11118 4917 11118 4 _090_
rlabel metal1 s 4503 11798 4503 11798 4 _091_
rlabel metal2 s 2162 11730 2162 11730 4 _092_
rlabel metal1 s 1748 11322 1748 11322 4 _093_
rlabel metal1 s 2238 9962 2238 9962 4 _094_
rlabel metal2 s 2254 9350 2254 9350 4 _095_
rlabel metal2 s 10350 12002 10350 12002 4 _096_
rlabel metal1 s 12558 14960 12558 14960 4 _097_
rlabel metal2 s 12650 14144 12650 14144 4 _098_
rlabel metal1 s 15032 16082 15032 16082 4 _099_
rlabel metal2 s 14398 18530 14398 18530 4 _100_
rlabel metal2 s 16601 17646 16601 17646 4 _101_
rlabel metal1 s 18124 18938 18124 18938 4 _102_
rlabel metal1 s 17300 21930 17300 21930 4 _103_
rlabel metal2 s 14306 21794 14306 21794 4 _104_
rlabel metal1 s 12220 13226 12220 13226 4 _105_
rlabel metal1 s 3404 13838 3404 13838 4 _106_
rlabel metal1 s 3174 14484 3174 14484 4 _107_
rlabel metal1 s 2157 15062 2157 15062 4 _108_
rlabel metal1 s 2300 16150 2300 16150 4 _109_
rlabel metal1 s 2295 17170 2295 17170 4 _110_
rlabel metal2 s 2806 18530 2806 18530 4 _111_
rlabel metal1 s 2295 19346 2295 19346 4 _112_
rlabel metal1 s 3031 21590 3031 21590 4 _113_
rlabel metal1 s 17158 3910 17158 3910 4 _114_
rlabel metal1 s 16468 3978 16468 3978 4 _115_
rlabel metal2 s 16698 4420 16698 4420 4 _116_
rlabel metal1 s 17480 6834 17480 6834 4 _117_
rlabel metal1 s 19588 6630 19588 6630 4 _118_
rlabel metal1 s 19320 6970 19320 6970 4 _119_
rlabel metal2 s 19412 15674 19412 15674 4 _120_
rlabel metal2 s 19826 15674 19826 15674 4 _121_
rlabel metal1 s 18814 15028 18814 15028 4 _122_
rlabel metal1 s 14214 11322 14214 11322 4 _123_
rlabel metal1 s 14950 10778 14950 10778 4 _124_
rlabel metal1 s 14444 11254 14444 11254 4 _125_
rlabel metal1 s 5474 11322 5474 11322 4 _126_
rlabel metal2 s 6762 11016 6762 11016 4 _127_
rlabel metal1 s 7866 10676 7866 10676 4 _128_
rlabel metal1 s 20516 11322 20516 11322 4 _129_
rlabel metal2 s 20654 10234 20654 10234 4 _130_
rlabel metal1 s 21068 11322 21068 11322 4 _131_
rlabel metal1 s 9338 3400 9338 3400 4 _132_
rlabel metal1 s 8050 3536 8050 3536 4 _133_
rlabel metal1 s 7314 5168 7314 5168 4 _134_
rlabel metal1 s 7084 5202 7084 5202 4 _135_
rlabel metal2 s 7406 6800 7406 6800 4 _136_
rlabel metal1 s 12834 7888 12834 7888 4 _137_
rlabel metal1 s 7048 7271 7048 7271 4 _138_
rlabel metal1 s 6762 7514 6762 7514 4 _139_
rlabel metal1 s 7682 7412 7682 7412 4 _140_
rlabel metal2 s 7682 8262 7682 8262 4 _141_
rlabel metal1 s 7130 7276 7130 7276 4 _142_
rlabel metal1 s 6578 6358 6578 6358 4 _143_
rlabel metal1 s 7452 4590 7452 4590 4 _144_
rlabel metal1 s 7590 4726 7590 4726 4 _145_
rlabel metal1 s 7268 3706 7268 3706 4 _146_
rlabel metal2 s 8142 3978 8142 3978 4 _147_
rlabel metal1 s 8556 3026 8556 3026 4 _148_
rlabel metal1 s 2530 20978 2530 20978 4 _149_
rlabel metal1 s 3956 20570 3956 20570 4 _150_
rlabel metal1 s 4002 18768 4002 18768 4 _151_
rlabel metal1 s 4554 17510 4554 17510 4 _152_
rlabel metal2 s 5290 16524 5290 16524 4 _153_
rlabel metal1 s 5658 14450 5658 14450 4 _154_
rlabel metal1 s 7820 14314 7820 14314 4 _155_
rlabel metal1 s 5152 14586 5152 14586 4 _156_
rlabel metal1 s 4968 15402 4968 15402 4 _157_
rlabel metal1 s 4876 15130 4876 15130 4 _158_
rlabel metal1 s 4738 15504 4738 15504 4 _159_
rlabel metal1 s 4646 15674 4646 15674 4 _160_
rlabel metal1 s 4278 17306 4278 17306 4 _161_
rlabel metal2 s 4186 18496 4186 18496 4 _162_
rlabel metal1 s 4600 18734 4600 18734 4 _163_
rlabel metal1 s 3956 18938 3956 18938 4 _164_
rlabel metal1 s 2530 21386 2530 21386 4 _165_
rlabel metal1 s 13662 22542 13662 22542 4 _166_
rlabel metal1 s 13386 21556 13386 21556 4 _167_
rlabel metal1 s 12972 19890 12972 19890 4 _168_
rlabel metal1 s 12926 19414 12926 19414 4 _169_
rlabel metal1 s 12742 18292 12742 18292 4 _170_
rlabel metal1 s 13110 16524 13110 16524 4 _171_
rlabel metal1 s 12466 16456 12466 16456 4 _172_
rlabel metal2 s 12834 16966 12834 16966 4 _173_
rlabel metal1 s 13340 16626 13340 16626 4 _174_
rlabel metal2 s 12926 16966 12926 16966 4 _175_
rlabel metal1 s 12650 17136 12650 17136 4 _176_
rlabel metal1 s 12512 17306 12512 17306 4 _177_
rlabel metal1 s 13248 18394 13248 18394 4 _178_
rlabel metal1 s 13386 19482 13386 19482 4 _179_
rlabel metal1 s 13064 19822 13064 19822 4 _180_
rlabel metal1 s 13616 20026 13616 20026 4 _181_
rlabel metal1 s 13340 21658 13340 21658 4 _182_
rlabel metal1 s 17158 3706 17158 3706 4 _183_
rlabel metal1 s 16008 3706 16008 3706 4 _184_
rlabel metal1 s 18170 6970 18170 6970 4 _185_
rlabel metal1 s 18078 7378 18078 7378 4 _186_
rlabel metal1 s 19090 14960 19090 14960 4 _187_
rlabel metal1 s 19366 14994 19366 14994 4 _188_
rlabel metal1 s 13248 10166 13248 10166 4 _189_
rlabel metal1 s 14720 11322 14720 11322 4 _190_
rlabel metal1 s 3634 11288 3634 11288 4 _191_
rlabel metal1 s 7084 10778 7084 10778 4 _192_
rlabel metal2 s 19274 11492 19274 11492 4 _193_
rlabel metal2 s 20746 10948 20746 10948 4 _194_
rlabel metal2 s 14030 20196 14030 20196 4 _195_
rlabel metal1 s 8786 15538 8786 15538 4 _196_
rlabel metal1 s 12558 16048 12558 16048 4 _197_
rlabel metal1 s 12052 17646 12052 17646 4 _198_
rlabel metal1 s 10994 17748 10994 17748 4 _199_
rlabel metal1 s 10626 18938 10626 18938 4 _200_
rlabel metal1 s 17342 21590 17342 21590 4 _201_
rlabel metal1 s 2346 15538 2346 15538 4 _202_
rlabel metal1 s 11730 17850 11730 17850 4 _203_
rlabel metal1 s 5198 13872 5198 13872 4 _204_
rlabel metal1 s 10534 19380 10534 19380 4 _205_
rlabel metal1 s 10212 18734 10212 18734 4 _206_
rlabel metal2 s 10810 20944 10810 20944 4 _207_
rlabel metal2 s 10442 20774 10442 20774 4 _208_
rlabel metal2 s 12006 21539 12006 21539 4 _209_
rlabel metal1 s 10626 21488 10626 21488 4 _210_
rlabel metal1 s 12098 20570 12098 20570 4 _211_
rlabel metal1 s 17618 2448 17618 2448 4 _212_
rlabel metal1 s 16284 3026 16284 3026 4 _213_
rlabel metal1 s 13570 4114 13570 4114 4 _214_
rlabel metal2 s 13570 2587 13570 2587 4 _215_
rlabel metal1 s 17204 2414 17204 2414 4 _216_
rlabel metal1 s 18722 2482 18722 2482 4 _217_
rlabel metal1 s 16790 4692 16790 4692 4 _218_
rlabel metal1 s 18630 3706 18630 3706 4 _219_
rlabel metal1 s 20194 3162 20194 3162 4 _220_
rlabel metal1 s 18860 9554 18860 9554 4 _221_
rlabel metal1 s 18032 12818 18032 12818 4 _222_
rlabel metal1 s 20240 8942 20240 8942 4 _223_
rlabel metal1 s 21298 9622 21298 9622 4 _224_
rlabel metal1 s 18906 11220 18906 11220 4 _225_
rlabel metal1 s 19228 13294 19228 13294 4 _226_
rlabel metal1 s 17664 12614 17664 12614 4 _227_
rlabel metal1 s 19550 13328 19550 13328 4 _228_
rlabel metal1 s 20516 19822 20516 19822 4 _229_
rlabel metal2 s 12650 7106 12650 7106 4 _230_
rlabel metal1 s 13892 6358 13892 6358 4 _231_
rlabel metal1 s 13018 5678 13018 5678 4 _232_
rlabel metal1 s 12581 5542 12581 5542 4 _233_
rlabel metal1 s 9338 4114 9338 4114 4 _234_
rlabel metal2 s 11914 6596 11914 6596 4 _235_
rlabel metal1 s 12650 3570 12650 3570 4 _236_
rlabel metal1 s 11960 6290 11960 6290 4 _237_
rlabel metal1 s 8878 6766 8878 6766 4 _238_
rlabel metal1 s 10488 8534 10488 8534 4 _239_
rlabel metal1 s 11684 8942 11684 8942 4 _240_
rlabel metal1 s 10576 8602 10576 8602 4 _241_
rlabel metal2 s 11822 9350 11822 9350 4 _242_
rlabel metal1 s 13018 6970 13018 6970 4 _243_
rlabel metal1 s 13202 7514 13202 7514 4 _244_
rlabel metal2 s 12098 8500 12098 8500 4 _245_
rlabel metal1 s 9338 9044 9338 9044 4 _246_
rlabel metal1 s 9476 8602 9476 8602 4 _247_
rlabel metal1 s 9430 8908 9430 8908 4 _248_
rlabel metal2 s 10166 8330 10166 8330 4 _249_
rlabel metal1 s 9246 9996 9246 9996 4 _250_
rlabel metal1 s 9982 9690 9982 9690 4 _251_
rlabel metal1 s 8970 8432 8970 8432 4 _252_
rlabel metal1 s 8464 9146 8464 9146 4 _253_
rlabel metal1 s 8418 8976 8418 8976 4 _254_
rlabel metal1 s 8694 6324 8694 6324 4 _255_
rlabel metal1 s 8924 8058 8924 8058 4 _256_
rlabel metal1 s 9476 6766 9476 6766 4 _257_
rlabel metal1 s 8602 6358 8602 6358 4 _258_
rlabel metal1 s 6302 17238 6302 17238 4 _259_
rlabel metal1 s 8418 6358 8418 6358 4 _260_
rlabel metal1 s 9982 6698 9982 6698 4 _261_
rlabel metal1 s 9890 5882 9890 5882 4 _262_
rlabel metal2 s 9246 6596 9246 6596 4 _263_
rlabel metal1 s 10074 6868 10074 6868 4 _264_
rlabel metal1 s 10258 6800 10258 6800 4 _265_
rlabel metal2 s 12466 3434 12466 3434 4 _266_
rlabel metal1 s 11178 2890 11178 2890 4 _267_
rlabel metal1 s 10258 5338 10258 5338 4 _268_
rlabel metal1 s 10672 3366 10672 3366 4 _269_
rlabel metal1 s 11132 3910 11132 3910 4 _270_
rlabel metal1 s 12788 3706 12788 3706 4 _271_
rlabel metal1 s 11546 4113 11546 4113 4 _272_
rlabel metal1 s 12098 3536 12098 3536 4 _273_
rlabel metal1 s 9798 3400 9798 3400 4 _274_
rlabel metal1 s 9660 3706 9660 3706 4 _275_
rlabel metal1 s 9844 4114 9844 4114 4 _276_
rlabel metal2 s 10718 3774 10718 3774 4 _277_
rlabel metal1 s 10166 3638 10166 3638 4 _278_
rlabel metal1 s 15548 6290 15548 6290 4 _279_
rlabel metal1 s 16284 12818 16284 12818 4 _280_
rlabel metal1 s 20194 7820 20194 7820 4 _281_
rlabel metal1 s 21390 5338 21390 5338 4 _282_
rlabel metal1 s 20470 14926 20470 14926 4 _283_
rlabel metal1 s 20516 5338 20516 5338 4 _284_
rlabel metal1 s 18860 6766 18860 6766 4 _285_
rlabel metal1 s 16468 8466 16468 8466 4 _286_
rlabel metal2 s 16698 7378 16698 7378 4 _287_
rlabel metal1 s 16008 5678 16008 5678 4 _288_
rlabel metal1 s 13524 3706 13524 3706 4 _289_
rlabel metal1 s 20700 14994 20700 14994 4 _290_
rlabel metal1 s 20010 16150 20010 16150 4 _291_
rlabel metal1 s 19780 16762 19780 16762 4 _292_
rlabel metal1 s 17710 16524 17710 16524 4 _293_
rlabel metal1 s 18446 15402 18446 15402 4 _294_
rlabel metal1 s 17066 13906 17066 13906 4 _295_
rlabel metal1 s 18308 14042 18308 14042 4 _296_
rlabel metal1 s 17802 13940 17802 13940 4 _297_
rlabel metal1 s 19228 19346 19228 19346 4 _298_
rlabel metal1 s 13938 7854 13938 7854 4 _299_
rlabel metal1 s 9384 13362 9384 13362 4 _300_
rlabel metal2 s 9338 13872 9338 13872 4 _301_
rlabel metal2 s 9430 13872 9430 13872 4 _302_
rlabel metal1 s 5382 16014 5382 16014 4 _303_
rlabel metal2 s 7498 13804 7498 13804 4 _304_
rlabel metal1 s 7682 14416 7682 14416 4 _305_
rlabel metal1 s 7084 14246 7084 14246 4 _306_
rlabel metal1 s 8280 13294 8280 13294 4 _307_
rlabel metal1 s 6716 18870 6716 18870 4 _308_
rlabel metal1 s 6302 14314 6302 14314 4 _309_
rlabel metal1 s 6486 13838 6486 13838 4 _310_
rlabel metal1 s 7222 12750 7222 12750 4 _311_
rlabel metal1 s 7406 12852 7406 12852 4 _312_
rlabel metal1 s 9246 13770 9246 13770 4 _313_
rlabel metal1 s 8970 13804 8970 13804 4 _314_
rlabel metal1 s 8510 13974 8510 13974 4 _315_
rlabel metal2 s 7498 16252 7498 16252 4 _316_
rlabel metal1 s 8096 17102 8096 17102 4 _317_
rlabel metal1 s 8004 17034 8004 17034 4 _318_
rlabel metal1 s 7544 15470 7544 15470 4 _319_
rlabel metal2 s 7314 16422 7314 16422 4 _320_
rlabel metal2 s 7866 16422 7866 16422 4 _321_
rlabel metal1 s 6670 16592 6670 16592 4 _322_
rlabel metal1 s 6624 15946 6624 15946 4 _323_
rlabel metal1 s 6026 16082 6026 16082 4 _324_
rlabel metal1 s 6670 19414 6670 19414 4 _325_
rlabel metal1 s 6854 16218 6854 16218 4 _326_
rlabel metal1 s 6348 18258 6348 18258 4 _327_
rlabel metal1 s 5980 18394 5980 18394 4 _328_
rlabel metal2 s 6578 18700 6578 18700 4 _329_
rlabel metal1 s 8234 19278 8234 19278 4 _330_
rlabel metal1 s 6578 18666 6578 18666 4 _331_
rlabel metal1 s 7176 18734 7176 18734 4 _332_
rlabel metal2 s 8326 18904 8326 18904 4 _333_
rlabel metal1 s 8694 19346 8694 19346 4 _334_
rlabel metal2 s 7406 21114 7406 21114 4 _335_
rlabel metal1 s 6808 21454 6808 21454 4 _336_
rlabel metal1 s 7590 18190 7590 18190 4 _337_
rlabel metal1 s 7268 18394 7268 18394 4 _338_
rlabel metal2 s 8464 21114 8464 21114 4 _339_
rlabel metal1 s 8359 20774 8359 20774 4 _340_
rlabel metal2 s 8326 21556 8326 21556 4 _341_
rlabel metal1 s 6853 21522 6853 21522 4 _342_
rlabel metal1 s 6992 21046 6992 21046 4 _343_
rlabel metal1 s 5658 21590 5658 21590 4 _344_
rlabel metal1 s 6210 21012 6210 21012 4 _345_
rlabel metal1 s 6578 21114 6578 21114 4 _346_
rlabel metal1 s 6118 21318 6118 21318 4 _347_
rlabel metal1 s 11270 14042 11270 14042 4 _348_
rlabel metal1 s 5474 9588 5474 9588 4 _349_
rlabel metal1 s 4002 6324 4002 6324 4 _350_
rlabel metal1 s 5980 9010 5980 9010 4 _351_
rlabel metal1 s 5842 6358 5842 6358 4 _352_
rlabel metal1 s 5106 6290 5106 6290 4 _353_
rlabel metal1 s 5566 4692 5566 4692 4 _354_
rlabel metal1 s 4738 5236 4738 5236 4 _355_
rlabel metal1 s 5704 4522 5704 4522 4 _356_
rlabel metal1 s 4876 4114 4876 4114 4 _357_
rlabel metal1 s 8096 4114 8096 4114 4 _358_
rlabel metal1 s 5612 3162 5612 3162 4 _359_
rlabel metal1 s 8556 3706 8556 3706 4 _360_
rlabel metal1 s 16422 10642 16422 10642 4 _361_
rlabel metal1 s 16836 9690 16836 9690 4 _362_
rlabel metal1 s 15226 10132 15226 10132 4 _363_
rlabel metal1 s 14076 9622 14076 9622 4 _364_
rlabel metal2 s 12558 10982 12558 10982 4 _365_
rlabel metal1 s 11454 10778 11454 10778 4 _366_
rlabel metal1 s 2438 11152 2438 11152 4 _367_
rlabel metal1 s 10350 11220 10350 11220 4 _368_
rlabel metal1 s 14858 7854 14858 7854 4 _369_
rlabel metal1 s 7544 10642 7544 10642 4 _370_
rlabel metal1 s 6072 12206 6072 12206 4 _371_
rlabel metal1 s 5152 10234 5152 10234 4 _372_
rlabel metal1 s 4186 12614 4186 12614 4 _373_
rlabel metal1 s 1978 11084 1978 11084 4 _374_
rlabel metal1 s 1886 11152 1886 11152 4 _375_
rlabel metal1 s 1932 10030 1932 10030 4 _376_
rlabel metal1 s 2300 8942 2300 8942 4 _377_
rlabel metal1 s 10396 11730 10396 11730 4 _378_
rlabel metal1 s 16422 14008 16422 14008 4 _379_
rlabel metal1 s 15456 13498 15456 13498 4 _380_
rlabel metal1 s 15088 14450 15088 14450 4 _381_
rlabel metal1 s 15824 14042 15824 14042 4 _382_
rlabel metal1 s 15410 17612 15410 17612 4 _383_
rlabel metal1 s 14858 21522 14858 21522 4 _384_
rlabel metal1 s 14950 13770 14950 13770 4 _385_
rlabel metal2 s 15410 16898 15410 16898 4 _386_
rlabel metal2 s 15778 20230 15778 20230 4 _387_
rlabel metal1 s 15870 20230 15870 20230 4 _388_
rlabel metal1 s 13156 15674 13156 15674 4 _389_
rlabel metal1 s 13424 15334 13424 15334 4 _390_
rlabel metal2 s 12834 15232 12834 15232 4 _391_
rlabel metal2 s 14582 14688 14582 14688 4 _392_
rlabel metal2 s 15226 14790 15226 14790 4 _393_
rlabel metal1 s 13938 14382 13938 14382 4 _394_
rlabel metal1 s 12834 14416 12834 14416 4 _395_
rlabel metal1 s 14766 17136 14766 17136 4 _396_
rlabel metal1 s 15088 17170 15088 17170 4 _397_
rlabel metal1 s 14674 17238 14674 17238 4 _398_
rlabel metal1 s 14812 16422 14812 16422 4 _399_
rlabel metal1 s 14122 16082 14122 16082 4 _400_
rlabel metal1 s 14720 15674 14720 15674 4 _401_
rlabel metal1 s 14991 18190 14991 18190 4 _402_
rlabel metal2 s 14766 17680 14766 17680 4 _403_
rlabel metal1 s 14628 18258 14628 18258 4 _404_
rlabel metal1 s 16698 18700 16698 18700 4 _405_
rlabel metal1 s 15042 17680 15042 17680 4 _406_
rlabel metal1 s 16054 17748 16054 17748 4 _407_
rlabel metal2 s 17066 17952 17066 17952 4 _408_
rlabel metal1 s 16882 18190 16882 18190 4 _409_
rlabel metal2 s 18170 19210 18170 19210 4 _410_
rlabel metal1 s 16646 19368 16646 19368 4 _411_
rlabel metal1 s 17112 19210 17112 19210 4 _412_
rlabel metal1 s 17342 18938 17342 18938 4 _413_
rlabel metal1 s 17710 18802 17710 18802 4 _414_
rlabel metal1 s 16606 21114 16606 21114 4 _415_
rlabel metal1 s 16146 21386 16146 21386 4 _416_
rlabel metal2 s 16974 19686 16974 19686 4 _417_
rlabel metal1 s 16330 20400 16330 20400 4 _418_
rlabel metal2 s 16698 20910 16698 20910 4 _419_
rlabel metal1 s 15824 21454 15824 21454 4 _420_
rlabel metal1 s 17434 21352 17434 21352 4 _421_
rlabel metal1 s 17283 21658 17283 21658 4 _422_
rlabel metal1 s 17066 21318 17066 21318 4 _423_
rlabel metal1 s 15686 21046 15686 21046 4 _424_
rlabel metal2 s 15594 20740 15594 20740 4 _425_
rlabel metal1 s 14950 21012 14950 21012 4 _426_
rlabel metal1 s 14444 21114 14444 21114 4 _427_
rlabel metal1 s 15226 21114 15226 21114 4 _428_
rlabel metal1 s 11546 12206 11546 12206 4 _429_
rlabel metal1 s 4741 14042 4741 14042 4 _430_
rlabel metal1 s 2438 15436 2438 15436 4 _431_
rlabel metal1 s 4830 14892 4830 14892 4 _432_
rlabel metal2 s 3266 16524 3266 16524 4 _433_
rlabel metal2 s 2346 15878 2346 15878 4 _434_
rlabel metal1 s 3404 17646 3404 17646 4 _435_
rlabel metal1 s 3312 17170 3312 17170 4 _436_
rlabel metal1 s 3082 19788 3082 19788 4 _437_
rlabel metal2 s 2990 18972 2990 18972 4 _438_
rlabel metal2 s 3450 21556 3450 21556 4 _439_
rlabel metal2 s 3082 19516 3082 19516 4 _440_
rlabel metal1 s 3174 21114 3174 21114 4 _441_
rlabel metal2 s 11730 15606 11730 15606 4 clk
rlabel metal1 s 16514 5270 16514 5270 4 clknet_0_clk
rlabel metal1 s 1564 11730 1564 11730 4 clknet_3_0__leaf_clk
rlabel metal2 s 5566 4862 5566 4862 4 clknet_3_1__leaf_clk
rlabel metal1 s 2714 21420 2714 21420 4 clknet_3_2__leaf_clk
rlabel metal2 s 12098 13600 12098 13600 4 clknet_3_3__leaf_clk
rlabel metal1 s 13202 3978 13202 3978 4 clknet_3_4__leaf_clk
rlabel metal2 s 20562 9248 20562 9248 4 clknet_3_5__leaf_clk
rlabel metal2 s 19366 18258 19366 18258 4 clknet_3_6__leaf_clk
rlabel metal1 s 20010 13940 20010 13940 4 clknet_3_7__leaf_clk
rlabel metal1 s 14628 6630 14628 6630 4 d0.debounced
rlabel metal1 s 16514 3468 16514 3468 4 d0.state\[0\]
rlabel metal1 s 15962 4148 15962 4148 4 d0.state\[1\]
rlabel metal1 s 14812 4046 14812 4046 4 d0.state\[2\]
rlabel metal2 s 16146 3876 16146 3876 4 d0.state\[3\]
rlabel metal1 s 18354 2822 18354 2822 4 d0.state\[4\]
rlabel metal1 s 18124 4250 18124 4250 4 d0.state\[5\]
rlabel metal1 s 18124 3910 18124 3910 4 d0.state\[6\]
rlabel metal2 s 17894 3383 17894 3383 4 d0.state\[7\]
rlabel metal1 s 16974 7446 16974 7446 4 d1.debounced
rlabel metal1 s 20286 7174 20286 7174 4 d1.state\[0\]
rlabel metal1 s 20470 7514 20470 7514 4 d1.state\[1\]
rlabel metal1 s 21114 6086 21114 6086 4 d1.state\[2\]
rlabel metal2 s 19918 7140 19918 7140 4 d1.state\[3\]
rlabel metal2 s 18078 8092 18078 8092 4 d1.state\[4\]
rlabel metal2 s 17710 8228 17710 8228 4 d1.state\[5\]
rlabel metal1 s 17848 6698 17848 6698 4 d1.state\[6\]
rlabel metal1 s 15686 6222 15686 6222 4 d1.state\[7\]
rlabel metal1 s 14490 13974 14490 13974 4 d3.debounced
rlabel metal1 s 21114 15674 21114 15674 4 d3.state\[0\]
rlabel metal2 s 21666 16388 21666 16388 4 d3.state\[1\]
rlabel metal1 s 21390 17306 21390 17306 4 d3.state\[2\]
rlabel metal1 s 20240 16626 20240 16626 4 d3.state\[3\]
rlabel metal2 s 18446 15130 18446 15130 4 d3.state\[4\]
rlabel metal1 s 17112 15470 17112 15470 4 d3.state\[5\]
rlabel metal1 s 18446 15062 18446 15062 4 d3.state\[6\]
rlabel metal1 s 18952 16626 18952 16626 4 d3.state\[7\]
rlabel metal1 s 13018 11662 13018 11662 4 d4.debounced
rlabel metal1 s 15640 11322 15640 11322 4 d4.state\[0\]
rlabel metal1 s 17112 10778 17112 10778 4 d4.state\[1\]
rlabel metal1 s 16882 10132 16882 10132 4 d4.state\[2\]
rlabel metal1 s 15180 11118 15180 11118 4 d4.state\[3\]
rlabel metal1 s 14030 10234 14030 10234 4 d4.state\[4\]
rlabel metal2 s 12650 10982 12650 10982 4 d4.state\[5\]
rlabel metal1 s 13478 11016 13478 11016 4 d4.state\[6\]
rlabel metal1 s 13432 10098 13432 10098 4 d4.state\[7\]
rlabel metal1 s 14306 13158 14306 13158 4 d5.debounced
rlabel metal1 s 6762 11254 6762 11254 4 d5.state\[0\]
rlabel metal1 s 6302 10778 6302 10778 4 d5.state\[1\]
rlabel metal2 s 6578 10302 6578 10302 4 d5.state\[2\]
rlabel metal1 s 5980 10098 5980 10098 4 d5.state\[3\]
rlabel metal1 s 3588 12342 3588 12342 4 d5.state\[4\]
rlabel metal1 s 3726 11628 3726 11628 4 d5.state\[5\]
rlabel metal1 s 3634 10642 3634 10642 4 d5.state\[6\]
rlabel metal1 s 3082 10574 3082 10574 4 d5.state\[7\]
rlabel metal1 s 15870 12716 15870 12716 4 d6.debounced
rlabel metal1 s 20608 10234 20608 10234 4 d6.state\[0\]
rlabel metal1 s 19136 9690 19136 9690 4 d6.state\[1\]
rlabel metal1 s 21160 9962 21160 9962 4 d6.state\[2\]
rlabel metal2 s 21022 9690 21022 9690 4 d6.state\[3\]
rlabel metal1 s 19780 11322 19780 11322 4 d6.state\[4\]
rlabel metal1 s 19412 12206 19412 12206 4 d6.state\[5\]
rlabel metal1 s 21068 12954 21068 12954 4 d6.state\[6\]
rlabel metal1 s 21482 13294 21482 13294 4 d6.state\[7\]
rlabel metal1 s 13662 6868 13662 6868 4 e0.old_a
rlabel metal1 s 15042 7310 15042 7310 4 e0.old_b
rlabel metal1 s 12788 7990 12788 7990 4 e0.value\[0\]
rlabel metal1 s 12834 8602 12834 8602 4 e0.value\[1\]
rlabel metal2 s 8418 8364 8418 8364 4 e0.value\[2\]
rlabel metal1 s 7406 8806 7406 8806 4 e0.value\[3\]
rlabel metal1 s 7682 6290 7682 6290 4 e0.value\[4\]
rlabel metal1 s 9430 6290 9430 6290 4 e0.value\[5\]
rlabel metal1 s 11546 3910 11546 3910 4 e0.value\[6\]
rlabel metal1 s 10764 3162 10764 3162 4 e0.value\[7\]
rlabel metal1 s 10120 14042 10120 14042 4 e1.old_a
rlabel metal1 s 10810 13362 10810 13362 4 e1.old_b
rlabel metal1 s 6900 13294 6900 13294 4 e1.value\[0\]
rlabel metal1 s 8510 14314 8510 14314 4 e1.value\[1\]
rlabel metal2 s 8602 16014 8602 16014 4 e1.value\[2\]
rlabel metal1 s 5842 16762 5842 16762 4 e1.value\[3\]
rlabel metal2 s 5566 17952 5566 17952 4 e1.value\[4\]
rlabel metal1 s 7912 18598 7912 18598 4 e1.value\[5\]
rlabel metal2 s 6670 21148 6670 21148 4 e1.value\[6\]
rlabel metal1 s 6854 21862 6854 21862 4 e1.value\[7\]
rlabel metal1 s 14076 13362 14076 13362 4 e2.old_a
rlabel metal2 s 15686 13600 15686 13600 4 e2.old_b
rlabel metal1 s 13202 15470 13202 15470 4 e2.value\[0\]
rlabel metal1 s 13202 16592 13202 16592 4 e2.value\[1\]
rlabel metal2 s 13478 17102 13478 17102 4 e2.value\[2\]
rlabel metal1 s 13846 18258 13846 18258 4 e2.value\[3\]
rlabel metal2 s 17434 18598 17434 18598 4 e2.value\[4\]
rlabel metal1 s 13570 19788 13570 19788 4 e2.value\[5\]
rlabel metal1 s 13294 22134 13294 22134 4 e2.value\[6\]
rlabel metal1 s 13708 21522 13708 21522 4 e2.value\[7\]
rlabel metal1 s 21942 2414 21942 2414 4 enc0_a
rlabel metal2 s 46 1588 46 1588 4 enc0_b
rlabel metal1 s 19504 22610 19504 22610 4 enc1_a
rlabel metal2 s 17434 823 17434 823 4 enc1_b
rlabel metal3 s 820 8908 820 8908 4 enc2_a
rlabel metal1 s 21942 21522 21942 21522 4 enc2_b
rlabel metal1 s 20838 3026 20838 3026 4 net1
rlabel metal1 s 12098 22610 12098 22610 4 net10
rlabel metal2 s 12374 21182 12374 21182 4 net11
rlabel metal1 s 3496 21862 3496 21862 4 net12
rlabel metal1 s 8280 3978 8280 3978 4 net13
rlabel metal2 s 4002 14416 4002 14416 4 net14
rlabel metal1 s 12650 17544 12650 17544 4 net15
rlabel metal1 s 3404 19346 3404 19346 4 net16
rlabel metal1 s 5934 4114 5934 4114 4 net17
rlabel metal1 s 4186 9520 4186 9520 4 net18
rlabel metal1 s 10902 21556 10902 21556 4 net19
rlabel metal1 s 4255 2278 4255 2278 4 net2
rlabel metal2 s 11546 18564 11546 18564 4 net20
rlabel metal1 s 3542 17102 3542 17102 4 net21
rlabel metal1 s 21666 10166 21666 10166 4 net22
rlabel metal1 s 5336 5134 5336 5134 4 net23
rlabel metal2 s 16974 6970 16974 6970 4 net24
rlabel metal1 s 4508 15062 4508 15062 4 net25
rlabel metal1 s 2622 15504 2622 15504 4 net26
rlabel metal1 s 10534 17306 10534 17306 4 net27
rlabel metal2 s 9890 16558 9890 16558 4 net28
rlabel metal1 s 10902 20366 10902 20366 4 net29
rlabel metal1 s 19412 22406 19412 22406 4 net3
rlabel metal1 s 3358 18190 3358 18190 4 net30
rlabel metal1 s 13294 17102 13294 17102 4 net31
rlabel metal1 s 11285 16150 11285 16150 4 net32
rlabel metal2 s 11822 11084 11822 11084 4 net33
rlabel metal1 s 14720 3502 14720 3502 4 net34
rlabel metal2 s 6394 9078 6394 9078 4 net35
rlabel metal1 s 4278 8976 4278 8976 4 net36
rlabel metal1 s 7084 13158 7084 13158 4 net37
rlabel metal1 s 7084 10642 7084 10642 4 net38
rlabel metal1 s 4922 4012 4922 4012 4 net39
rlabel metal1 s 19136 2618 19136 2618 4 net4
rlabel metal1 s 13156 8942 13156 8942 4 net40
rlabel metal1 s 4002 14586 4002 14586 4 net41
rlabel metal2 s 18446 7242 18446 7242 4 net42
rlabel metal1 s 20010 5202 20010 5202 4 net43
rlabel metal1 s 20378 11866 20378 11866 4 net44
rlabel metal1 s 3082 10778 3082 10778 4 net45
rlabel metal1 s 3082 11254 3082 11254 4 net46
rlabel metal2 s 18446 9724 18446 9724 4 net47
rlabel metal1 s 21344 7922 21344 7922 4 net48
rlabel metal1 s 17894 2414 17894 2414 4 net49
rlabel metal1 s 1978 8976 1978 8976 4 net5
rlabel metal1 s 16054 10676 16054 10676 4 net50
rlabel metal1 s 20286 15062 20286 15062 4 net51
rlabel metal1 s 13754 9486 13754 9486 4 net52
rlabel metal1 s 3680 12410 3680 12410 4 net53
rlabel metal2 s 19090 16388 19090 16388 4 net54
rlabel metal2 s 11914 18496 11914 18496 4 net55
rlabel metal1 s 18032 5202 18032 5202 4 net56
rlabel metal1 s 20424 8602 20424 8602 4 net57
rlabel metal1 s 16422 11662 16422 11662 4 net58
rlabel metal2 s 5566 12036 5566 12036 4 net59
rlabel metal1 s 20516 20434 20516 20434 4 net6
rlabel metal1 s 16514 5814 16514 5814 4 net60
rlabel metal1 s 20930 16694 20930 16694 4 net61
rlabel metal1 s 5796 9146 5796 9146 4 net62
rlabel metal1 s 20976 13294 20976 13294 4 net63
rlabel metal1 s 18998 12342 18998 12342 4 net64
rlabel metal1 s 2576 10574 2576 10574 4 net65
rlabel metal1 s 12144 10098 12144 10098 4 net66
rlabel metal1 s 19642 15572 19642 15572 4 net67
rlabel metal1 s 18998 12818 18998 12818 4 net68
rlabel metal1 s 19182 3502 19182 3502 4 net69
rlabel metal1 s 15870 11798 15870 11798 4 net7
rlabel metal1 s 19596 16626 19596 16626 4 net70
rlabel metal1 s 17802 8602 17802 8602 4 net71
rlabel metal1 s 14260 4046 14260 4046 4 net72
rlabel metal2 s 20654 5372 20654 5372 4 net73
rlabel metal1 s 17480 3570 17480 3570 4 net74
rlabel metal2 s 12834 11186 12834 11186 4 net75
rlabel metal1 s 2530 15538 2530 15538 4 net76
rlabel metal2 s 15226 4454 15226 4454 4 net77
rlabel metal1 s 17296 9486 17296 9486 4 net78
rlabel metal1 s 17526 13838 17526 13838 4 net79
rlabel metal1 s 8832 2414 8832 2414 4 net8
rlabel metal1 s 4140 6290 4140 6290 4 net80
rlabel metal1 s 14030 15470 14030 15470 4 net81
rlabel metal1 s 5428 10030 5428 10030 4 net82
rlabel metal1 s 10718 3026 10718 3026 4 net83
rlabel metal1 s 6670 20468 6670 20468 4 net84
rlabel metal1 s 16606 14518 16606 14518 4 net85
rlabel metal2 s 11408 8602 11408 8602 4 net86
rlabel metal1 s 2070 21386 2070 21386 4 net9
rlabel metal2 s 6946 7548 6946 7548 4 p0.counter\[0\]
rlabel metal1 s 6072 8942 6072 8942 4 p0.counter\[1\]
rlabel metal1 s 5382 7174 5382 7174 4 p0.counter\[2\]
rlabel metal1 s 6762 6324 6762 6324 4 p0.counter\[3\]
rlabel metal1 s 5796 5678 5796 5678 4 p0.counter\[4\]
rlabel metal2 s 7682 4675 7682 4675 4 p0.counter\[5\]
rlabel metal1 s 7222 3638 7222 3638 4 p0.counter\[6\]
rlabel metal1 s 7130 4114 7130 4114 4 p0.counter\[7\]
rlabel metal1 s 4370 14382 4370 14382 4 p1.counter\[0\]
rlabel metal1 s 3404 14586 3404 14586 4 p1.counter\[1\]
rlabel metal2 s 4278 14977 4278 14977 4 p1.counter\[2\]
rlabel metal1 s 4646 16558 4646 16558 4 p1.counter\[3\]
rlabel metal1 s 4508 17714 4508 17714 4 p1.counter\[4\]
rlabel metal1 s 4646 18190 4646 18190 4 p1.counter\[5\]
rlabel metal1 s 3818 19448 3818 19448 4 p1.counter\[6\]
rlabel metal1 s 2622 21590 2622 21590 4 p1.counter\[7\]
rlabel metal1 s 10258 16966 10258 16966 4 p2.counter\[0\]
rlabel metal1 s 11960 17102 11960 17102 4 p2.counter\[1\]
rlabel metal2 s 11270 16898 11270 16898 4 p2.counter\[2\]
rlabel metal1 s 11960 18938 11960 18938 4 p2.counter\[3\]
rlabel metal2 s 12650 19006 12650 19006 4 p2.counter\[4\]
rlabel metal1 s 12466 20468 12466 20468 4 p2.counter\[5\]
rlabel metal1 s 12742 21012 12742 21012 4 p2.counter\[6\]
rlabel metal2 s 13110 21828 13110 21828 4 p2.counter\[7\]
rlabel metal2 s 8418 1520 8418 1520 4 pwm0_out
rlabel metal1 s 1426 22746 1426 22746 4 pwm1_out
rlabel metal1 s 10534 22746 10534 22746 4 pwm2_out
rlabel metal1 s 21666 11696 21666 11696 4 reset
flabel metal5 s 1056 20764 22312 21084 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 15596 22312 15916 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 10428 22312 10748 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 5260 22312 5580 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 20119 2128 20439 22896 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 14829 2128 15149 22896 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 9539 2128 9859 22896 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4249 2128 4569 22896 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 20104 22312 20424 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 14936 22312 15256 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 9768 22312 10088 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 4600 22312 4920 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 19459 2128 19779 22896 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 14169 2128 14489 22896 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 8879 2128 9199 22896 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3589 2128 3909 22896 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 18368 800 18488 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 22608 2048 23408 2168 0 FreeSans 600 0 0 0 enc0_a
port 4 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 enc0_b
port 5 nsew
flabel metal2 s 19338 24752 19394 25552 0 FreeSans 280 90 0 0 enc1_a
port 6 nsew
flabel metal2 s 17406 0 17462 800 0 FreeSans 280 90 0 0 enc1_b
port 7 nsew
flabel metal3 s 0 8848 800 8968 0 FreeSans 600 0 0 0 enc2_a
port 8 nsew
flabel metal3 s 22608 21088 23408 21208 0 FreeSans 600 0 0 0 enc2_b
port 9 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 pwm0_out
port 10 nsew
flabel metal2 s 1306 24752 1362 25552 0 FreeSans 280 90 0 0 pwm1_out
port 11 nsew
flabel metal2 s 10322 24752 10378 25552 0 FreeSans 280 90 0 0 pwm2_out
port 12 nsew
flabel metal3 s 22608 11568 23408 11688 0 FreeSans 600 0 0 0 reset
port 13 nsew
<< properties >>
string FIXED_BBOX 0 0 23408 25552
<< end >>
